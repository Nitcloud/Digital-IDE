.INIT_RAM_00({INIT[255:0]}),
.INIT_RAM_01({INIT[511:256]}),
.INIT_RAM_02({INIT[767:512]}),
.INIT_RAM_03({INIT[1023:768]}),
.INIT_RAM_04({INIT[1279:1024]}),
.INIT_RAM_05({INIT[1535:1280]}),
.INIT_RAM_06({INIT[1791:1536]}),
.INIT_RAM_07({INIT[2047:1792]}),
.INIT_RAM_08({INIT[2303:2048]}),
.INIT_RAM_09({INIT[2559:2304]}),
.INIT_RAM_0A({INIT[2815:2560]}),
.INIT_RAM_0B({INIT[3071:2816]}),
.INIT_RAM_0C({INIT[3327:3072]}),
.INIT_RAM_0D({INIT[3583:3328]}),
.INIT_RAM_0E({INIT[3839:3584]}),
.INIT_RAM_0F({INIT[4095:3840]}),
.INIT_RAM_10({INIT[4351:4096]}),
.INIT_RAM_11({INIT[4607:4352]}),
.INIT_RAM_12({INIT[4863:4608]}),
.INIT_RAM_13({INIT[5119:4864]}),
.INIT_RAM_14({INIT[5375:5120]}),
.INIT_RAM_15({INIT[5631:5376]}),
.INIT_RAM_16({INIT[5887:5632]}),
.INIT_RAM_17({INIT[6143:5888]}),
.INIT_RAM_18({INIT[6399:6144]}),
.INIT_RAM_19({INIT[6655:6400]}),
.INIT_RAM_1A({INIT[6911:6656]}),
.INIT_RAM_1B({INIT[7167:6912]}),
.INIT_RAM_1C({INIT[7423:7168]}),
.INIT_RAM_1D({INIT[7679:7424]}),
.INIT_RAM_1E({INIT[7935:7680]}),
.INIT_RAM_1F({INIT[8191:7936]}),
.INIT_RAM_20({INIT[8447:8192]}),
.INIT_RAM_21({INIT[8703:8448]}),
.INIT_RAM_22({INIT[8959:8704]}),
.INIT_RAM_23({INIT[9215:8960]}),
.INIT_RAM_24({INIT[9471:9216]}),
.INIT_RAM_25({INIT[9727:9472]}),
.INIT_RAM_26({INIT[9983:9728]}),
.INIT_RAM_27({INIT[10239:9984]}),
.INIT_RAM_28({INIT[10495:10240]}),
.INIT_RAM_29({INIT[10751:10496]}),
.INIT_RAM_2A({INIT[11007:10752]}),
.INIT_RAM_2B({INIT[11263:11008]}),
.INIT_RAM_2C({INIT[11519:11264]}),
.INIT_RAM_2D({INIT[11775:11520]}),
.INIT_RAM_2E({INIT[12031:11776]}),
.INIT_RAM_2F({INIT[12287:12032]}),
.INIT_RAM_30({INIT[12543:12288]}),
.INIT_RAM_31({INIT[12799:12544]}),
.INIT_RAM_32({INIT[13055:12800]}),
.INIT_RAM_33({INIT[13311:13056]}),
.INIT_RAM_34({INIT[13567:13312]}),
.INIT_RAM_35({INIT[13823:13568]}),
.INIT_RAM_36({INIT[14079:13824]}),
.INIT_RAM_37({INIT[14335:14080]}),
.INIT_RAM_38({INIT[14591:14336]}),
.INIT_RAM_39({INIT[14847:14592]}),
.INIT_RAM_3A({INIT[15103:14848]}),
.INIT_RAM_3B({INIT[15359:15104]}),
.INIT_RAM_3C({INIT[15615:15360]}),
.INIT_RAM_3D({INIT[15871:15616]}),
.INIT_RAM_3E({INIT[16127:15872]}),
.INIT_RAM_3F({INIT[16383:16128]}),
