.INIT_00(INIT[  0*256 +: 256]),
.INIT_01(INIT[  1*256 +: 256]),
.INIT_02(INIT[  2*256 +: 256]),
.INIT_03(INIT[  3*256 +: 256]),
.INIT_04(INIT[  4*256 +: 256]),
.INIT_05(INIT[  5*256 +: 256]),
.INIT_06(INIT[  6*256 +: 256]),
.INIT_07(INIT[  7*256 +: 256]),
.INIT_08(INIT[  8*256 +: 256]),
.INIT_09(INIT[  9*256 +: 256]),
.INIT_0A(INIT[ 10*256 +: 256]),
.INIT_0B(INIT[ 11*256 +: 256]),
.INIT_0C(INIT[ 12*256 +: 256]),
.INIT_0D(INIT[ 13*256 +: 256]),
.INIT_0E(INIT[ 14*256 +: 256]),
.INIT_0F(INIT[ 15*256 +: 256]),
.INIT_10(INIT[ 16*256 +: 256]),
.INIT_11(INIT[ 17*256 +: 256]),
.INIT_12(INIT[ 18*256 +: 256]),
.INIT_13(INIT[ 19*256 +: 256]),
.INIT_14(INIT[ 20*256 +: 256]),
.INIT_15(INIT[ 21*256 +: 256]),
.INIT_16(INIT[ 22*256 +: 256]),
.INIT_17(INIT[ 23*256 +: 256]),
.INIT_18(INIT[ 24*256 +: 256]),
.INIT_19(INIT[ 25*256 +: 256]),
.INIT_1A(INIT[ 26*256 +: 256]),
.INIT_1B(INIT[ 27*256 +: 256]),
.INIT_1C(INIT[ 28*256 +: 256]),
.INIT_1D(INIT[ 29*256 +: 256]),
.INIT_1E(INIT[ 30*256 +: 256]),
.INIT_1F(INIT[ 31*256 +: 256]),
