    .ADA0(1'b0), .ADA1(1'b0), .ADA2(A1ADDR[0]), .ADA3(A1ADDR[1]), .ADA4(A1ADDR[2]), .ADA5(A1ADDR[3]), .ADA6(A1ADDR[4]), .ADA7(A1ADDR[5]), .ADA8(A1ADDR[6]), .ADA9(A1ADDR[7]), .ADA10(A1ADDR[8]), .ADA11(A1ADDR[9]), .ADA12(A1ADDR[10]), .ADA13(A1ADDR[11]),
    .ADB0(1'b0), .ADB1(1'b0), .ADB2(B1ADDR[0]), .ADB3(B1ADDR[1]), .ADB4(B1ADDR[2]), .ADB5(B1ADDR[3]), .ADB6(B1ADDR[4]), .ADB7(B1ADDR[5]), .ADB8(B1ADDR[6]), .ADB9(B1ADDR[7]), .ADB10(B1ADDR[8]), .ADB11(B1ADDR[9]), .ADB12(B1ADDR[10]), .ADB13(B1ADDR[11]),
    .DIA0(A1DATA[0]), .DIA1(A1DATA[1]), .DIA2(A1DATA[2]), .DIA3(A1DATA[3]), .DIA4(1'b0), .DIA5(1'b0), .DIA6(1'b0), .DIA7(1'b0), .DIA8(1'b0), .DIA9(1'b0), .DIA10(1'b0), .DIA11(1'b0), .DIA12(1'b0), .DIA13(1'b0), .DIA14(1'b0), .DIA15(1'b0), .DIA16(1'b0), .DIA17(1'b0),
    .DOB0(B1DATA[0]), .DOB1(B1DATA[1]), .DOB2(B1DATA[2]), .DOB3(B1DATA[3]),
