.INITP_00({ INIT[255*9+8], INIT[254*9+8], INIT[253*9+8], INIT[252*9+8],
            INIT[251*9+8], INIT[250*9+8], INIT[249*9+8], INIT[248*9+8],
            INIT[247*9+8], INIT[246*9+8], INIT[245*9+8], INIT[244*9+8],
            INIT[243*9+8], INIT[242*9+8], INIT[241*9+8], INIT[240*9+8],
            INIT[239*9+8], INIT[238*9+8], INIT[237*9+8], INIT[236*9+8],
            INIT[235*9+8], INIT[234*9+8], INIT[233*9+8], INIT[232*9+8],
            INIT[231*9+8], INIT[230*9+8], INIT[229*9+8], INIT[228*9+8],
            INIT[227*9+8], INIT[226*9+8], INIT[225*9+8], INIT[224*9+8],
            INIT[223*9+8], INIT[222*9+8], INIT[221*9+8], INIT[220*9+8],
            INIT[219*9+8], INIT[218*9+8], INIT[217*9+8], INIT[216*9+8],
            INIT[215*9+8], INIT[214*9+8], INIT[213*9+8], INIT[212*9+8],
            INIT[211*9+8], INIT[210*9+8], INIT[209*9+8], INIT[208*9+8],
            INIT[207*9+8], INIT[206*9+8], INIT[205*9+8], INIT[204*9+8],
            INIT[203*9+8], INIT[202*9+8], INIT[201*9+8], INIT[200*9+8],
            INIT[199*9+8], INIT[198*9+8], INIT[197*9+8], INIT[196*9+8],
            INIT[195*9+8], INIT[194*9+8], INIT[193*9+8], INIT[192*9+8],
            INIT[191*9+8], INIT[190*9+8], INIT[189*9+8], INIT[188*9+8],
            INIT[187*9+8], INIT[186*9+8], INIT[185*9+8], INIT[184*9+8],
            INIT[183*9+8], INIT[182*9+8], INIT[181*9+8], INIT[180*9+8],
            INIT[179*9+8], INIT[178*9+8], INIT[177*9+8], INIT[176*9+8],
            INIT[175*9+8], INIT[174*9+8], INIT[173*9+8], INIT[172*9+8],
            INIT[171*9+8], INIT[170*9+8], INIT[169*9+8], INIT[168*9+8],
            INIT[167*9+8], INIT[166*9+8], INIT[165*9+8], INIT[164*9+8],
            INIT[163*9+8], INIT[162*9+8], INIT[161*9+8], INIT[160*9+8],
            INIT[159*9+8], INIT[158*9+8], INIT[157*9+8], INIT[156*9+8],
            INIT[155*9+8], INIT[154*9+8], INIT[153*9+8], INIT[152*9+8],
            INIT[151*9+8], INIT[150*9+8], INIT[149*9+8], INIT[148*9+8],
            INIT[147*9+8], INIT[146*9+8], INIT[145*9+8], INIT[144*9+8],
            INIT[143*9+8], INIT[142*9+8], INIT[141*9+8], INIT[140*9+8],
            INIT[139*9+8], INIT[138*9+8], INIT[137*9+8], INIT[136*9+8],
            INIT[135*9+8], INIT[134*9+8], INIT[133*9+8], INIT[132*9+8],
            INIT[131*9+8], INIT[130*9+8], INIT[129*9+8], INIT[128*9+8],
            INIT[127*9+8], INIT[126*9+8], INIT[125*9+8], INIT[124*9+8],
            INIT[123*9+8], INIT[122*9+8], INIT[121*9+8], INIT[120*9+8],
            INIT[119*9+8], INIT[118*9+8], INIT[117*9+8], INIT[116*9+8],
            INIT[115*9+8], INIT[114*9+8], INIT[113*9+8], INIT[112*9+8],
            INIT[111*9+8], INIT[110*9+8], INIT[109*9+8], INIT[108*9+8],
            INIT[107*9+8], INIT[106*9+8], INIT[105*9+8], INIT[104*9+8],
            INIT[103*9+8], INIT[102*9+8], INIT[101*9+8], INIT[100*9+8],
            INIT[ 99*9+8], INIT[ 98*9+8], INIT[ 97*9+8], INIT[ 96*9+8],
            INIT[ 95*9+8], INIT[ 94*9+8], INIT[ 93*9+8], INIT[ 92*9+8],
            INIT[ 91*9+8], INIT[ 90*9+8], INIT[ 89*9+8], INIT[ 88*9+8],
            INIT[ 87*9+8], INIT[ 86*9+8], INIT[ 85*9+8], INIT[ 84*9+8],
            INIT[ 83*9+8], INIT[ 82*9+8], INIT[ 81*9+8], INIT[ 80*9+8],
            INIT[ 79*9+8], INIT[ 78*9+8], INIT[ 77*9+8], INIT[ 76*9+8],
            INIT[ 75*9+8], INIT[ 74*9+8], INIT[ 73*9+8], INIT[ 72*9+8],
            INIT[ 71*9+8], INIT[ 70*9+8], INIT[ 69*9+8], INIT[ 68*9+8],
            INIT[ 67*9+8], INIT[ 66*9+8], INIT[ 65*9+8], INIT[ 64*9+8],
            INIT[ 63*9+8], INIT[ 62*9+8], INIT[ 61*9+8], INIT[ 60*9+8],
            INIT[ 59*9+8], INIT[ 58*9+8], INIT[ 57*9+8], INIT[ 56*9+8],
            INIT[ 55*9+8], INIT[ 54*9+8], INIT[ 53*9+8], INIT[ 52*9+8],
            INIT[ 51*9+8], INIT[ 50*9+8], INIT[ 49*9+8], INIT[ 48*9+8],
            INIT[ 47*9+8], INIT[ 46*9+8], INIT[ 45*9+8], INIT[ 44*9+8],
            INIT[ 43*9+8], INIT[ 42*9+8], INIT[ 41*9+8], INIT[ 40*9+8],
            INIT[ 39*9+8], INIT[ 38*9+8], INIT[ 37*9+8], INIT[ 36*9+8],
            INIT[ 35*9+8], INIT[ 34*9+8], INIT[ 33*9+8], INIT[ 32*9+8],
            INIT[ 31*9+8], INIT[ 30*9+8], INIT[ 29*9+8], INIT[ 28*9+8],
            INIT[ 27*9+8], INIT[ 26*9+8], INIT[ 25*9+8], INIT[ 24*9+8],
            INIT[ 23*9+8], INIT[ 22*9+8], INIT[ 21*9+8], INIT[ 20*9+8],
            INIT[ 19*9+8], INIT[ 18*9+8], INIT[ 17*9+8], INIT[ 16*9+8],
            INIT[ 15*9+8], INIT[ 14*9+8], INIT[ 13*9+8], INIT[ 12*9+8],
            INIT[ 11*9+8], INIT[ 10*9+8], INIT[  9*9+8], INIT[  8*9+8],
            INIT[  7*9+8], INIT[  6*9+8], INIT[  5*9+8], INIT[  4*9+8],
            INIT[  3*9+8], INIT[  2*9+8], INIT[  1*9+8], INIT[  0*9+8]}),
.INITP_01({ INIT[511*9+8], INIT[510*9+8], INIT[509*9+8], INIT[508*9+8],
            INIT[507*9+8], INIT[506*9+8], INIT[505*9+8], INIT[504*9+8],
            INIT[503*9+8], INIT[502*9+8], INIT[501*9+8], INIT[500*9+8],
            INIT[499*9+8], INIT[498*9+8], INIT[497*9+8], INIT[496*9+8],
            INIT[495*9+8], INIT[494*9+8], INIT[493*9+8], INIT[492*9+8],
            INIT[491*9+8], INIT[490*9+8], INIT[489*9+8], INIT[488*9+8],
            INIT[487*9+8], INIT[486*9+8], INIT[485*9+8], INIT[484*9+8],
            INIT[483*9+8], INIT[482*9+8], INIT[481*9+8], INIT[480*9+8],
            INIT[479*9+8], INIT[478*9+8], INIT[477*9+8], INIT[476*9+8],
            INIT[475*9+8], INIT[474*9+8], INIT[473*9+8], INIT[472*9+8],
            INIT[471*9+8], INIT[470*9+8], INIT[469*9+8], INIT[468*9+8],
            INIT[467*9+8], INIT[466*9+8], INIT[465*9+8], INIT[464*9+8],
            INIT[463*9+8], INIT[462*9+8], INIT[461*9+8], INIT[460*9+8],
            INIT[459*9+8], INIT[458*9+8], INIT[457*9+8], INIT[456*9+8],
            INIT[455*9+8], INIT[454*9+8], INIT[453*9+8], INIT[452*9+8],
            INIT[451*9+8], INIT[450*9+8], INIT[449*9+8], INIT[448*9+8],
            INIT[447*9+8], INIT[446*9+8], INIT[445*9+8], INIT[444*9+8],
            INIT[443*9+8], INIT[442*9+8], INIT[441*9+8], INIT[440*9+8],
            INIT[439*9+8], INIT[438*9+8], INIT[437*9+8], INIT[436*9+8],
            INIT[435*9+8], INIT[434*9+8], INIT[433*9+8], INIT[432*9+8],
            INIT[431*9+8], INIT[430*9+8], INIT[429*9+8], INIT[428*9+8],
            INIT[427*9+8], INIT[426*9+8], INIT[425*9+8], INIT[424*9+8],
            INIT[423*9+8], INIT[422*9+8], INIT[421*9+8], INIT[420*9+8],
            INIT[419*9+8], INIT[418*9+8], INIT[417*9+8], INIT[416*9+8],
            INIT[415*9+8], INIT[414*9+8], INIT[413*9+8], INIT[412*9+8],
            INIT[411*9+8], INIT[410*9+8], INIT[409*9+8], INIT[408*9+8],
            INIT[407*9+8], INIT[406*9+8], INIT[405*9+8], INIT[404*9+8],
            INIT[403*9+8], INIT[402*9+8], INIT[401*9+8], INIT[400*9+8],
            INIT[399*9+8], INIT[398*9+8], INIT[397*9+8], INIT[396*9+8],
            INIT[395*9+8], INIT[394*9+8], INIT[393*9+8], INIT[392*9+8],
            INIT[391*9+8], INIT[390*9+8], INIT[389*9+8], INIT[388*9+8],
            INIT[387*9+8], INIT[386*9+8], INIT[385*9+8], INIT[384*9+8],
            INIT[383*9+8], INIT[382*9+8], INIT[381*9+8], INIT[380*9+8],
            INIT[379*9+8], INIT[378*9+8], INIT[377*9+8], INIT[376*9+8],
            INIT[375*9+8], INIT[374*9+8], INIT[373*9+8], INIT[372*9+8],
            INIT[371*9+8], INIT[370*9+8], INIT[369*9+8], INIT[368*9+8],
            INIT[367*9+8], INIT[366*9+8], INIT[365*9+8], INIT[364*9+8],
            INIT[363*9+8], INIT[362*9+8], INIT[361*9+8], INIT[360*9+8],
            INIT[359*9+8], INIT[358*9+8], INIT[357*9+8], INIT[356*9+8],
            INIT[355*9+8], INIT[354*9+8], INIT[353*9+8], INIT[352*9+8],
            INIT[351*9+8], INIT[350*9+8], INIT[349*9+8], INIT[348*9+8],
            INIT[347*9+8], INIT[346*9+8], INIT[345*9+8], INIT[344*9+8],
            INIT[343*9+8], INIT[342*9+8], INIT[341*9+8], INIT[340*9+8],
            INIT[339*9+8], INIT[338*9+8], INIT[337*9+8], INIT[336*9+8],
            INIT[335*9+8], INIT[334*9+8], INIT[333*9+8], INIT[332*9+8],
            INIT[331*9+8], INIT[330*9+8], INIT[329*9+8], INIT[328*9+8],
            INIT[327*9+8], INIT[326*9+8], INIT[325*9+8], INIT[324*9+8],
            INIT[323*9+8], INIT[322*9+8], INIT[321*9+8], INIT[320*9+8],
            INIT[319*9+8], INIT[318*9+8], INIT[317*9+8], INIT[316*9+8],
            INIT[315*9+8], INIT[314*9+8], INIT[313*9+8], INIT[312*9+8],
            INIT[311*9+8], INIT[310*9+8], INIT[309*9+8], INIT[308*9+8],
            INIT[307*9+8], INIT[306*9+8], INIT[305*9+8], INIT[304*9+8],
            INIT[303*9+8], INIT[302*9+8], INIT[301*9+8], INIT[300*9+8],
            INIT[299*9+8], INIT[298*9+8], INIT[297*9+8], INIT[296*9+8],
            INIT[295*9+8], INIT[294*9+8], INIT[293*9+8], INIT[292*9+8],
            INIT[291*9+8], INIT[290*9+8], INIT[289*9+8], INIT[288*9+8],
            INIT[287*9+8], INIT[286*9+8], INIT[285*9+8], INIT[284*9+8],
            INIT[283*9+8], INIT[282*9+8], INIT[281*9+8], INIT[280*9+8],
            INIT[279*9+8], INIT[278*9+8], INIT[277*9+8], INIT[276*9+8],
            INIT[275*9+8], INIT[274*9+8], INIT[273*9+8], INIT[272*9+8],
            INIT[271*9+8], INIT[270*9+8], INIT[269*9+8], INIT[268*9+8],
            INIT[267*9+8], INIT[266*9+8], INIT[265*9+8], INIT[264*9+8],
            INIT[263*9+8], INIT[262*9+8], INIT[261*9+8], INIT[260*9+8],
            INIT[259*9+8], INIT[258*9+8], INIT[257*9+8], INIT[256*9+8]}),
.INITP_02({ INIT[767*9+8], INIT[766*9+8], INIT[765*9+8], INIT[764*9+8],
            INIT[763*9+8], INIT[762*9+8], INIT[761*9+8], INIT[760*9+8],
            INIT[759*9+8], INIT[758*9+8], INIT[757*9+8], INIT[756*9+8],
            INIT[755*9+8], INIT[754*9+8], INIT[753*9+8], INIT[752*9+8],
            INIT[751*9+8], INIT[750*9+8], INIT[749*9+8], INIT[748*9+8],
            INIT[747*9+8], INIT[746*9+8], INIT[745*9+8], INIT[744*9+8],
            INIT[743*9+8], INIT[742*9+8], INIT[741*9+8], INIT[740*9+8],
            INIT[739*9+8], INIT[738*9+8], INIT[737*9+8], INIT[736*9+8],
            INIT[735*9+8], INIT[734*9+8], INIT[733*9+8], INIT[732*9+8],
            INIT[731*9+8], INIT[730*9+8], INIT[729*9+8], INIT[728*9+8],
            INIT[727*9+8], INIT[726*9+8], INIT[725*9+8], INIT[724*9+8],
            INIT[723*9+8], INIT[722*9+8], INIT[721*9+8], INIT[720*9+8],
            INIT[719*9+8], INIT[718*9+8], INIT[717*9+8], INIT[716*9+8],
            INIT[715*9+8], INIT[714*9+8], INIT[713*9+8], INIT[712*9+8],
            INIT[711*9+8], INIT[710*9+8], INIT[709*9+8], INIT[708*9+8],
            INIT[707*9+8], INIT[706*9+8], INIT[705*9+8], INIT[704*9+8],
            INIT[703*9+8], INIT[702*9+8], INIT[701*9+8], INIT[700*9+8],
            INIT[699*9+8], INIT[698*9+8], INIT[697*9+8], INIT[696*9+8],
            INIT[695*9+8], INIT[694*9+8], INIT[693*9+8], INIT[692*9+8],
            INIT[691*9+8], INIT[690*9+8], INIT[689*9+8], INIT[688*9+8],
            INIT[687*9+8], INIT[686*9+8], INIT[685*9+8], INIT[684*9+8],
            INIT[683*9+8], INIT[682*9+8], INIT[681*9+8], INIT[680*9+8],
            INIT[679*9+8], INIT[678*9+8], INIT[677*9+8], INIT[676*9+8],
            INIT[675*9+8], INIT[674*9+8], INIT[673*9+8], INIT[672*9+8],
            INIT[671*9+8], INIT[670*9+8], INIT[669*9+8], INIT[668*9+8],
            INIT[667*9+8], INIT[666*9+8], INIT[665*9+8], INIT[664*9+8],
            INIT[663*9+8], INIT[662*9+8], INIT[661*9+8], INIT[660*9+8],
            INIT[659*9+8], INIT[658*9+8], INIT[657*9+8], INIT[656*9+8],
            INIT[655*9+8], INIT[654*9+8], INIT[653*9+8], INIT[652*9+8],
            INIT[651*9+8], INIT[650*9+8], INIT[649*9+8], INIT[648*9+8],
            INIT[647*9+8], INIT[646*9+8], INIT[645*9+8], INIT[644*9+8],
            INIT[643*9+8], INIT[642*9+8], INIT[641*9+8], INIT[640*9+8],
            INIT[639*9+8], INIT[638*9+8], INIT[637*9+8], INIT[636*9+8],
            INIT[635*9+8], INIT[634*9+8], INIT[633*9+8], INIT[632*9+8],
            INIT[631*9+8], INIT[630*9+8], INIT[629*9+8], INIT[628*9+8],
            INIT[627*9+8], INIT[626*9+8], INIT[625*9+8], INIT[624*9+8],
            INIT[623*9+8], INIT[622*9+8], INIT[621*9+8], INIT[620*9+8],
            INIT[619*9+8], INIT[618*9+8], INIT[617*9+8], INIT[616*9+8],
            INIT[615*9+8], INIT[614*9+8], INIT[613*9+8], INIT[612*9+8],
            INIT[611*9+8], INIT[610*9+8], INIT[609*9+8], INIT[608*9+8],
            INIT[607*9+8], INIT[606*9+8], INIT[605*9+8], INIT[604*9+8],
            INIT[603*9+8], INIT[602*9+8], INIT[601*9+8], INIT[600*9+8],
            INIT[599*9+8], INIT[598*9+8], INIT[597*9+8], INIT[596*9+8],
            INIT[595*9+8], INIT[594*9+8], INIT[593*9+8], INIT[592*9+8],
            INIT[591*9+8], INIT[590*9+8], INIT[589*9+8], INIT[588*9+8],
            INIT[587*9+8], INIT[586*9+8], INIT[585*9+8], INIT[584*9+8],
            INIT[583*9+8], INIT[582*9+8], INIT[581*9+8], INIT[580*9+8],
            INIT[579*9+8], INIT[578*9+8], INIT[577*9+8], INIT[576*9+8],
            INIT[575*9+8], INIT[574*9+8], INIT[573*9+8], INIT[572*9+8],
            INIT[571*9+8], INIT[570*9+8], INIT[569*9+8], INIT[568*9+8],
            INIT[567*9+8], INIT[566*9+8], INIT[565*9+8], INIT[564*9+8],
            INIT[563*9+8], INIT[562*9+8], INIT[561*9+8], INIT[560*9+8],
            INIT[559*9+8], INIT[558*9+8], INIT[557*9+8], INIT[556*9+8],
            INIT[555*9+8], INIT[554*9+8], INIT[553*9+8], INIT[552*9+8],
            INIT[551*9+8], INIT[550*9+8], INIT[549*9+8], INIT[548*9+8],
            INIT[547*9+8], INIT[546*9+8], INIT[545*9+8], INIT[544*9+8],
            INIT[543*9+8], INIT[542*9+8], INIT[541*9+8], INIT[540*9+8],
            INIT[539*9+8], INIT[538*9+8], INIT[537*9+8], INIT[536*9+8],
            INIT[535*9+8], INIT[534*9+8], INIT[533*9+8], INIT[532*9+8],
            INIT[531*9+8], INIT[530*9+8], INIT[529*9+8], INIT[528*9+8],
            INIT[527*9+8], INIT[526*9+8], INIT[525*9+8], INIT[524*9+8],
            INIT[523*9+8], INIT[522*9+8], INIT[521*9+8], INIT[520*9+8],
            INIT[519*9+8], INIT[518*9+8], INIT[517*9+8], INIT[516*9+8],
            INIT[515*9+8], INIT[514*9+8], INIT[513*9+8], INIT[512*9+8]}),
.INITP_03({ INIT[1023*9+8], INIT[1022*9+8], INIT[1021*9+8], INIT[1020*9+8],
            INIT[1019*9+8], INIT[1018*9+8], INIT[1017*9+8], INIT[1016*9+8],
            INIT[1015*9+8], INIT[1014*9+8], INIT[1013*9+8], INIT[1012*9+8],
            INIT[1011*9+8], INIT[1010*9+8], INIT[1009*9+8], INIT[1008*9+8],
            INIT[1007*9+8], INIT[1006*9+8], INIT[1005*9+8], INIT[1004*9+8],
            INIT[1003*9+8], INIT[1002*9+8], INIT[1001*9+8], INIT[1000*9+8],
            INIT[999*9+8], INIT[998*9+8], INIT[997*9+8], INIT[996*9+8],
            INIT[995*9+8], INIT[994*9+8], INIT[993*9+8], INIT[992*9+8],
            INIT[991*9+8], INIT[990*9+8], INIT[989*9+8], INIT[988*9+8],
            INIT[987*9+8], INIT[986*9+8], INIT[985*9+8], INIT[984*9+8],
            INIT[983*9+8], INIT[982*9+8], INIT[981*9+8], INIT[980*9+8],
            INIT[979*9+8], INIT[978*9+8], INIT[977*9+8], INIT[976*9+8],
            INIT[975*9+8], INIT[974*9+8], INIT[973*9+8], INIT[972*9+8],
            INIT[971*9+8], INIT[970*9+8], INIT[969*9+8], INIT[968*9+8],
            INIT[967*9+8], INIT[966*9+8], INIT[965*9+8], INIT[964*9+8],
            INIT[963*9+8], INIT[962*9+8], INIT[961*9+8], INIT[960*9+8],
            INIT[959*9+8], INIT[958*9+8], INIT[957*9+8], INIT[956*9+8],
            INIT[955*9+8], INIT[954*9+8], INIT[953*9+8], INIT[952*9+8],
            INIT[951*9+8], INIT[950*9+8], INIT[949*9+8], INIT[948*9+8],
            INIT[947*9+8], INIT[946*9+8], INIT[945*9+8], INIT[944*9+8],
            INIT[943*9+8], INIT[942*9+8], INIT[941*9+8], INIT[940*9+8],
            INIT[939*9+8], INIT[938*9+8], INIT[937*9+8], INIT[936*9+8],
            INIT[935*9+8], INIT[934*9+8], INIT[933*9+8], INIT[932*9+8],
            INIT[931*9+8], INIT[930*9+8], INIT[929*9+8], INIT[928*9+8],
            INIT[927*9+8], INIT[926*9+8], INIT[925*9+8], INIT[924*9+8],
            INIT[923*9+8], INIT[922*9+8], INIT[921*9+8], INIT[920*9+8],
            INIT[919*9+8], INIT[918*9+8], INIT[917*9+8], INIT[916*9+8],
            INIT[915*9+8], INIT[914*9+8], INIT[913*9+8], INIT[912*9+8],
            INIT[911*9+8], INIT[910*9+8], INIT[909*9+8], INIT[908*9+8],
            INIT[907*9+8], INIT[906*9+8], INIT[905*9+8], INIT[904*9+8],
            INIT[903*9+8], INIT[902*9+8], INIT[901*9+8], INIT[900*9+8],
            INIT[899*9+8], INIT[898*9+8], INIT[897*9+8], INIT[896*9+8],
            INIT[895*9+8], INIT[894*9+8], INIT[893*9+8], INIT[892*9+8],
            INIT[891*9+8], INIT[890*9+8], INIT[889*9+8], INIT[888*9+8],
            INIT[887*9+8], INIT[886*9+8], INIT[885*9+8], INIT[884*9+8],
            INIT[883*9+8], INIT[882*9+8], INIT[881*9+8], INIT[880*9+8],
            INIT[879*9+8], INIT[878*9+8], INIT[877*9+8], INIT[876*9+8],
            INIT[875*9+8], INIT[874*9+8], INIT[873*9+8], INIT[872*9+8],
            INIT[871*9+8], INIT[870*9+8], INIT[869*9+8], INIT[868*9+8],
            INIT[867*9+8], INIT[866*9+8], INIT[865*9+8], INIT[864*9+8],
            INIT[863*9+8], INIT[862*9+8], INIT[861*9+8], INIT[860*9+8],
            INIT[859*9+8], INIT[858*9+8], INIT[857*9+8], INIT[856*9+8],
            INIT[855*9+8], INIT[854*9+8], INIT[853*9+8], INIT[852*9+8],
            INIT[851*9+8], INIT[850*9+8], INIT[849*9+8], INIT[848*9+8],
            INIT[847*9+8], INIT[846*9+8], INIT[845*9+8], INIT[844*9+8],
            INIT[843*9+8], INIT[842*9+8], INIT[841*9+8], INIT[840*9+8],
            INIT[839*9+8], INIT[838*9+8], INIT[837*9+8], INIT[836*9+8],
            INIT[835*9+8], INIT[834*9+8], INIT[833*9+8], INIT[832*9+8],
            INIT[831*9+8], INIT[830*9+8], INIT[829*9+8], INIT[828*9+8],
            INIT[827*9+8], INIT[826*9+8], INIT[825*9+8], INIT[824*9+8],
            INIT[823*9+8], INIT[822*9+8], INIT[821*9+8], INIT[820*9+8],
            INIT[819*9+8], INIT[818*9+8], INIT[817*9+8], INIT[816*9+8],
            INIT[815*9+8], INIT[814*9+8], INIT[813*9+8], INIT[812*9+8],
            INIT[811*9+8], INIT[810*9+8], INIT[809*9+8], INIT[808*9+8],
            INIT[807*9+8], INIT[806*9+8], INIT[805*9+8], INIT[804*9+8],
            INIT[803*9+8], INIT[802*9+8], INIT[801*9+8], INIT[800*9+8],
            INIT[799*9+8], INIT[798*9+8], INIT[797*9+8], INIT[796*9+8],
            INIT[795*9+8], INIT[794*9+8], INIT[793*9+8], INIT[792*9+8],
            INIT[791*9+8], INIT[790*9+8], INIT[789*9+8], INIT[788*9+8],
            INIT[787*9+8], INIT[786*9+8], INIT[785*9+8], INIT[784*9+8],
            INIT[783*9+8], INIT[782*9+8], INIT[781*9+8], INIT[780*9+8],
            INIT[779*9+8], INIT[778*9+8], INIT[777*9+8], INIT[776*9+8],
            INIT[775*9+8], INIT[774*9+8], INIT[773*9+8], INIT[772*9+8],
            INIT[771*9+8], INIT[770*9+8], INIT[769*9+8], INIT[768*9+8]}),
.INIT_00({ INIT[ 31*9 +: 8], INIT[ 30*9 +: 8], INIT[ 29*9 +: 8], INIT[ 28*9 +: 8],
           INIT[ 27*9 +: 8], INIT[ 26*9 +: 8], INIT[ 25*9 +: 8], INIT[ 24*9 +: 8],
           INIT[ 23*9 +: 8], INIT[ 22*9 +: 8], INIT[ 21*9 +: 8], INIT[ 20*9 +: 8],
           INIT[ 19*9 +: 8], INIT[ 18*9 +: 8], INIT[ 17*9 +: 8], INIT[ 16*9 +: 8],
           INIT[ 15*9 +: 8], INIT[ 14*9 +: 8], INIT[ 13*9 +: 8], INIT[ 12*9 +: 8],
           INIT[ 11*9 +: 8], INIT[ 10*9 +: 8], INIT[  9*9 +: 8], INIT[  8*9 +: 8],
           INIT[  7*9 +: 8], INIT[  6*9 +: 8], INIT[  5*9 +: 8], INIT[  4*9 +: 8],
           INIT[  3*9 +: 8], INIT[  2*9 +: 8], INIT[  1*9 +: 8], INIT[  0*9 +: 8]}),
.INIT_01({ INIT[ 63*9 +: 8], INIT[ 62*9 +: 8], INIT[ 61*9 +: 8], INIT[ 60*9 +: 8],
           INIT[ 59*9 +: 8], INIT[ 58*9 +: 8], INIT[ 57*9 +: 8], INIT[ 56*9 +: 8],
           INIT[ 55*9 +: 8], INIT[ 54*9 +: 8], INIT[ 53*9 +: 8], INIT[ 52*9 +: 8],
           INIT[ 51*9 +: 8], INIT[ 50*9 +: 8], INIT[ 49*9 +: 8], INIT[ 48*9 +: 8],
           INIT[ 47*9 +: 8], INIT[ 46*9 +: 8], INIT[ 45*9 +: 8], INIT[ 44*9 +: 8],
           INIT[ 43*9 +: 8], INIT[ 42*9 +: 8], INIT[ 41*9 +: 8], INIT[ 40*9 +: 8],
           INIT[ 39*9 +: 8], INIT[ 38*9 +: 8], INIT[ 37*9 +: 8], INIT[ 36*9 +: 8],
           INIT[ 35*9 +: 8], INIT[ 34*9 +: 8], INIT[ 33*9 +: 8], INIT[ 32*9 +: 8]}),
.INIT_02({ INIT[ 95*9 +: 8], INIT[ 94*9 +: 8], INIT[ 93*9 +: 8], INIT[ 92*9 +: 8],
           INIT[ 91*9 +: 8], INIT[ 90*9 +: 8], INIT[ 89*9 +: 8], INIT[ 88*9 +: 8],
           INIT[ 87*9 +: 8], INIT[ 86*9 +: 8], INIT[ 85*9 +: 8], INIT[ 84*9 +: 8],
           INIT[ 83*9 +: 8], INIT[ 82*9 +: 8], INIT[ 81*9 +: 8], INIT[ 80*9 +: 8],
           INIT[ 79*9 +: 8], INIT[ 78*9 +: 8], INIT[ 77*9 +: 8], INIT[ 76*9 +: 8],
           INIT[ 75*9 +: 8], INIT[ 74*9 +: 8], INIT[ 73*9 +: 8], INIT[ 72*9 +: 8],
           INIT[ 71*9 +: 8], INIT[ 70*9 +: 8], INIT[ 69*9 +: 8], INIT[ 68*9 +: 8],
           INIT[ 67*9 +: 8], INIT[ 66*9 +: 8], INIT[ 65*9 +: 8], INIT[ 64*9 +: 8]}),
.INIT_03({ INIT[127*9 +: 8], INIT[126*9 +: 8], INIT[125*9 +: 8], INIT[124*9 +: 8],
           INIT[123*9 +: 8], INIT[122*9 +: 8], INIT[121*9 +: 8], INIT[120*9 +: 8],
           INIT[119*9 +: 8], INIT[118*9 +: 8], INIT[117*9 +: 8], INIT[116*9 +: 8],
           INIT[115*9 +: 8], INIT[114*9 +: 8], INIT[113*9 +: 8], INIT[112*9 +: 8],
           INIT[111*9 +: 8], INIT[110*9 +: 8], INIT[109*9 +: 8], INIT[108*9 +: 8],
           INIT[107*9 +: 8], INIT[106*9 +: 8], INIT[105*9 +: 8], INIT[104*9 +: 8],
           INIT[103*9 +: 8], INIT[102*9 +: 8], INIT[101*9 +: 8], INIT[100*9 +: 8],
           INIT[ 99*9 +: 8], INIT[ 98*9 +: 8], INIT[ 97*9 +: 8], INIT[ 96*9 +: 8]}),
.INIT_04({ INIT[159*9 +: 8], INIT[158*9 +: 8], INIT[157*9 +: 8], INIT[156*9 +: 8],
           INIT[155*9 +: 8], INIT[154*9 +: 8], INIT[153*9 +: 8], INIT[152*9 +: 8],
           INIT[151*9 +: 8], INIT[150*9 +: 8], INIT[149*9 +: 8], INIT[148*9 +: 8],
           INIT[147*9 +: 8], INIT[146*9 +: 8], INIT[145*9 +: 8], INIT[144*9 +: 8],
           INIT[143*9 +: 8], INIT[142*9 +: 8], INIT[141*9 +: 8], INIT[140*9 +: 8],
           INIT[139*9 +: 8], INIT[138*9 +: 8], INIT[137*9 +: 8], INIT[136*9 +: 8],
           INIT[135*9 +: 8], INIT[134*9 +: 8], INIT[133*9 +: 8], INIT[132*9 +: 8],
           INIT[131*9 +: 8], INIT[130*9 +: 8], INIT[129*9 +: 8], INIT[128*9 +: 8]}),
.INIT_05({ INIT[191*9 +: 8], INIT[190*9 +: 8], INIT[189*9 +: 8], INIT[188*9 +: 8],
           INIT[187*9 +: 8], INIT[186*9 +: 8], INIT[185*9 +: 8], INIT[184*9 +: 8],
           INIT[183*9 +: 8], INIT[182*9 +: 8], INIT[181*9 +: 8], INIT[180*9 +: 8],
           INIT[179*9 +: 8], INIT[178*9 +: 8], INIT[177*9 +: 8], INIT[176*9 +: 8],
           INIT[175*9 +: 8], INIT[174*9 +: 8], INIT[173*9 +: 8], INIT[172*9 +: 8],
           INIT[171*9 +: 8], INIT[170*9 +: 8], INIT[169*9 +: 8], INIT[168*9 +: 8],
           INIT[167*9 +: 8], INIT[166*9 +: 8], INIT[165*9 +: 8], INIT[164*9 +: 8],
           INIT[163*9 +: 8], INIT[162*9 +: 8], INIT[161*9 +: 8], INIT[160*9 +: 8]}),
.INIT_06({ INIT[223*9 +: 8], INIT[222*9 +: 8], INIT[221*9 +: 8], INIT[220*9 +: 8],
           INIT[219*9 +: 8], INIT[218*9 +: 8], INIT[217*9 +: 8], INIT[216*9 +: 8],
           INIT[215*9 +: 8], INIT[214*9 +: 8], INIT[213*9 +: 8], INIT[212*9 +: 8],
           INIT[211*9 +: 8], INIT[210*9 +: 8], INIT[209*9 +: 8], INIT[208*9 +: 8],
           INIT[207*9 +: 8], INIT[206*9 +: 8], INIT[205*9 +: 8], INIT[204*9 +: 8],
           INIT[203*9 +: 8], INIT[202*9 +: 8], INIT[201*9 +: 8], INIT[200*9 +: 8],
           INIT[199*9 +: 8], INIT[198*9 +: 8], INIT[197*9 +: 8], INIT[196*9 +: 8],
           INIT[195*9 +: 8], INIT[194*9 +: 8], INIT[193*9 +: 8], INIT[192*9 +: 8]}),
.INIT_07({ INIT[255*9 +: 8], INIT[254*9 +: 8], INIT[253*9 +: 8], INIT[252*9 +: 8],
           INIT[251*9 +: 8], INIT[250*9 +: 8], INIT[249*9 +: 8], INIT[248*9 +: 8],
           INIT[247*9 +: 8], INIT[246*9 +: 8], INIT[245*9 +: 8], INIT[244*9 +: 8],
           INIT[243*9 +: 8], INIT[242*9 +: 8], INIT[241*9 +: 8], INIT[240*9 +: 8],
           INIT[239*9 +: 8], INIT[238*9 +: 8], INIT[237*9 +: 8], INIT[236*9 +: 8],
           INIT[235*9 +: 8], INIT[234*9 +: 8], INIT[233*9 +: 8], INIT[232*9 +: 8],
           INIT[231*9 +: 8], INIT[230*9 +: 8], INIT[229*9 +: 8], INIT[228*9 +: 8],
           INIT[227*9 +: 8], INIT[226*9 +: 8], INIT[225*9 +: 8], INIT[224*9 +: 8]}),
.INIT_08({ INIT[287*9 +: 8], INIT[286*9 +: 8], INIT[285*9 +: 8], INIT[284*9 +: 8],
           INIT[283*9 +: 8], INIT[282*9 +: 8], INIT[281*9 +: 8], INIT[280*9 +: 8],
           INIT[279*9 +: 8], INIT[278*9 +: 8], INIT[277*9 +: 8], INIT[276*9 +: 8],
           INIT[275*9 +: 8], INIT[274*9 +: 8], INIT[273*9 +: 8], INIT[272*9 +: 8],
           INIT[271*9 +: 8], INIT[270*9 +: 8], INIT[269*9 +: 8], INIT[268*9 +: 8],
           INIT[267*9 +: 8], INIT[266*9 +: 8], INIT[265*9 +: 8], INIT[264*9 +: 8],
           INIT[263*9 +: 8], INIT[262*9 +: 8], INIT[261*9 +: 8], INIT[260*9 +: 8],
           INIT[259*9 +: 8], INIT[258*9 +: 8], INIT[257*9 +: 8], INIT[256*9 +: 8]}),
.INIT_09({ INIT[319*9 +: 8], INIT[318*9 +: 8], INIT[317*9 +: 8], INIT[316*9 +: 8],
           INIT[315*9 +: 8], INIT[314*9 +: 8], INIT[313*9 +: 8], INIT[312*9 +: 8],
           INIT[311*9 +: 8], INIT[310*9 +: 8], INIT[309*9 +: 8], INIT[308*9 +: 8],
           INIT[307*9 +: 8], INIT[306*9 +: 8], INIT[305*9 +: 8], INIT[304*9 +: 8],
           INIT[303*9 +: 8], INIT[302*9 +: 8], INIT[301*9 +: 8], INIT[300*9 +: 8],
           INIT[299*9 +: 8], INIT[298*9 +: 8], INIT[297*9 +: 8], INIT[296*9 +: 8],
           INIT[295*9 +: 8], INIT[294*9 +: 8], INIT[293*9 +: 8], INIT[292*9 +: 8],
           INIT[291*9 +: 8], INIT[290*9 +: 8], INIT[289*9 +: 8], INIT[288*9 +: 8]}),
.INIT_0A({ INIT[351*9 +: 8], INIT[350*9 +: 8], INIT[349*9 +: 8], INIT[348*9 +: 8],
           INIT[347*9 +: 8], INIT[346*9 +: 8], INIT[345*9 +: 8], INIT[344*9 +: 8],
           INIT[343*9 +: 8], INIT[342*9 +: 8], INIT[341*9 +: 8], INIT[340*9 +: 8],
           INIT[339*9 +: 8], INIT[338*9 +: 8], INIT[337*9 +: 8], INIT[336*9 +: 8],
           INIT[335*9 +: 8], INIT[334*9 +: 8], INIT[333*9 +: 8], INIT[332*9 +: 8],
           INIT[331*9 +: 8], INIT[330*9 +: 8], INIT[329*9 +: 8], INIT[328*9 +: 8],
           INIT[327*9 +: 8], INIT[326*9 +: 8], INIT[325*9 +: 8], INIT[324*9 +: 8],
           INIT[323*9 +: 8], INIT[322*9 +: 8], INIT[321*9 +: 8], INIT[320*9 +: 8]}),
.INIT_0B({ INIT[383*9 +: 8], INIT[382*9 +: 8], INIT[381*9 +: 8], INIT[380*9 +: 8],
           INIT[379*9 +: 8], INIT[378*9 +: 8], INIT[377*9 +: 8], INIT[376*9 +: 8],
           INIT[375*9 +: 8], INIT[374*9 +: 8], INIT[373*9 +: 8], INIT[372*9 +: 8],
           INIT[371*9 +: 8], INIT[370*9 +: 8], INIT[369*9 +: 8], INIT[368*9 +: 8],
           INIT[367*9 +: 8], INIT[366*9 +: 8], INIT[365*9 +: 8], INIT[364*9 +: 8],
           INIT[363*9 +: 8], INIT[362*9 +: 8], INIT[361*9 +: 8], INIT[360*9 +: 8],
           INIT[359*9 +: 8], INIT[358*9 +: 8], INIT[357*9 +: 8], INIT[356*9 +: 8],
           INIT[355*9 +: 8], INIT[354*9 +: 8], INIT[353*9 +: 8], INIT[352*9 +: 8]}),
.INIT_0C({ INIT[415*9 +: 8], INIT[414*9 +: 8], INIT[413*9 +: 8], INIT[412*9 +: 8],
           INIT[411*9 +: 8], INIT[410*9 +: 8], INIT[409*9 +: 8], INIT[408*9 +: 8],
           INIT[407*9 +: 8], INIT[406*9 +: 8], INIT[405*9 +: 8], INIT[404*9 +: 8],
           INIT[403*9 +: 8], INIT[402*9 +: 8], INIT[401*9 +: 8], INIT[400*9 +: 8],
           INIT[399*9 +: 8], INIT[398*9 +: 8], INIT[397*9 +: 8], INIT[396*9 +: 8],
           INIT[395*9 +: 8], INIT[394*9 +: 8], INIT[393*9 +: 8], INIT[392*9 +: 8],
           INIT[391*9 +: 8], INIT[390*9 +: 8], INIT[389*9 +: 8], INIT[388*9 +: 8],
           INIT[387*9 +: 8], INIT[386*9 +: 8], INIT[385*9 +: 8], INIT[384*9 +: 8]}),
.INIT_0D({ INIT[447*9 +: 8], INIT[446*9 +: 8], INIT[445*9 +: 8], INIT[444*9 +: 8],
           INIT[443*9 +: 8], INIT[442*9 +: 8], INIT[441*9 +: 8], INIT[440*9 +: 8],
           INIT[439*9 +: 8], INIT[438*9 +: 8], INIT[437*9 +: 8], INIT[436*9 +: 8],
           INIT[435*9 +: 8], INIT[434*9 +: 8], INIT[433*9 +: 8], INIT[432*9 +: 8],
           INIT[431*9 +: 8], INIT[430*9 +: 8], INIT[429*9 +: 8], INIT[428*9 +: 8],
           INIT[427*9 +: 8], INIT[426*9 +: 8], INIT[425*9 +: 8], INIT[424*9 +: 8],
           INIT[423*9 +: 8], INIT[422*9 +: 8], INIT[421*9 +: 8], INIT[420*9 +: 8],
           INIT[419*9 +: 8], INIT[418*9 +: 8], INIT[417*9 +: 8], INIT[416*9 +: 8]}),
.INIT_0E({ INIT[479*9 +: 8], INIT[478*9 +: 8], INIT[477*9 +: 8], INIT[476*9 +: 8],
           INIT[475*9 +: 8], INIT[474*9 +: 8], INIT[473*9 +: 8], INIT[472*9 +: 8],
           INIT[471*9 +: 8], INIT[470*9 +: 8], INIT[469*9 +: 8], INIT[468*9 +: 8],
           INIT[467*9 +: 8], INIT[466*9 +: 8], INIT[465*9 +: 8], INIT[464*9 +: 8],
           INIT[463*9 +: 8], INIT[462*9 +: 8], INIT[461*9 +: 8], INIT[460*9 +: 8],
           INIT[459*9 +: 8], INIT[458*9 +: 8], INIT[457*9 +: 8], INIT[456*9 +: 8],
           INIT[455*9 +: 8], INIT[454*9 +: 8], INIT[453*9 +: 8], INIT[452*9 +: 8],
           INIT[451*9 +: 8], INIT[450*9 +: 8], INIT[449*9 +: 8], INIT[448*9 +: 8]}),
.INIT_0F({ INIT[511*9 +: 8], INIT[510*9 +: 8], INIT[509*9 +: 8], INIT[508*9 +: 8],
           INIT[507*9 +: 8], INIT[506*9 +: 8], INIT[505*9 +: 8], INIT[504*9 +: 8],
           INIT[503*9 +: 8], INIT[502*9 +: 8], INIT[501*9 +: 8], INIT[500*9 +: 8],
           INIT[499*9 +: 8], INIT[498*9 +: 8], INIT[497*9 +: 8], INIT[496*9 +: 8],
           INIT[495*9 +: 8], INIT[494*9 +: 8], INIT[493*9 +: 8], INIT[492*9 +: 8],
           INIT[491*9 +: 8], INIT[490*9 +: 8], INIT[489*9 +: 8], INIT[488*9 +: 8],
           INIT[487*9 +: 8], INIT[486*9 +: 8], INIT[485*9 +: 8], INIT[484*9 +: 8],
           INIT[483*9 +: 8], INIT[482*9 +: 8], INIT[481*9 +: 8], INIT[480*9 +: 8]}),
.INIT_10({ INIT[543*9 +: 8], INIT[542*9 +: 8], INIT[541*9 +: 8], INIT[540*9 +: 8],
           INIT[539*9 +: 8], INIT[538*9 +: 8], INIT[537*9 +: 8], INIT[536*9 +: 8],
           INIT[535*9 +: 8], INIT[534*9 +: 8], INIT[533*9 +: 8], INIT[532*9 +: 8],
           INIT[531*9 +: 8], INIT[530*9 +: 8], INIT[529*9 +: 8], INIT[528*9 +: 8],
           INIT[527*9 +: 8], INIT[526*9 +: 8], INIT[525*9 +: 8], INIT[524*9 +: 8],
           INIT[523*9 +: 8], INIT[522*9 +: 8], INIT[521*9 +: 8], INIT[520*9 +: 8],
           INIT[519*9 +: 8], INIT[518*9 +: 8], INIT[517*9 +: 8], INIT[516*9 +: 8],
           INIT[515*9 +: 8], INIT[514*9 +: 8], INIT[513*9 +: 8], INIT[512*9 +: 8]}),
.INIT_11({ INIT[575*9 +: 8], INIT[574*9 +: 8], INIT[573*9 +: 8], INIT[572*9 +: 8],
           INIT[571*9 +: 8], INIT[570*9 +: 8], INIT[569*9 +: 8], INIT[568*9 +: 8],
           INIT[567*9 +: 8], INIT[566*9 +: 8], INIT[565*9 +: 8], INIT[564*9 +: 8],
           INIT[563*9 +: 8], INIT[562*9 +: 8], INIT[561*9 +: 8], INIT[560*9 +: 8],
           INIT[559*9 +: 8], INIT[558*9 +: 8], INIT[557*9 +: 8], INIT[556*9 +: 8],
           INIT[555*9 +: 8], INIT[554*9 +: 8], INIT[553*9 +: 8], INIT[552*9 +: 8],
           INIT[551*9 +: 8], INIT[550*9 +: 8], INIT[549*9 +: 8], INIT[548*9 +: 8],
           INIT[547*9 +: 8], INIT[546*9 +: 8], INIT[545*9 +: 8], INIT[544*9 +: 8]}),
.INIT_12({ INIT[607*9 +: 8], INIT[606*9 +: 8], INIT[605*9 +: 8], INIT[604*9 +: 8],
           INIT[603*9 +: 8], INIT[602*9 +: 8], INIT[601*9 +: 8], INIT[600*9 +: 8],
           INIT[599*9 +: 8], INIT[598*9 +: 8], INIT[597*9 +: 8], INIT[596*9 +: 8],
           INIT[595*9 +: 8], INIT[594*9 +: 8], INIT[593*9 +: 8], INIT[592*9 +: 8],
           INIT[591*9 +: 8], INIT[590*9 +: 8], INIT[589*9 +: 8], INIT[588*9 +: 8],
           INIT[587*9 +: 8], INIT[586*9 +: 8], INIT[585*9 +: 8], INIT[584*9 +: 8],
           INIT[583*9 +: 8], INIT[582*9 +: 8], INIT[581*9 +: 8], INIT[580*9 +: 8],
           INIT[579*9 +: 8], INIT[578*9 +: 8], INIT[577*9 +: 8], INIT[576*9 +: 8]}),
.INIT_13({ INIT[639*9 +: 8], INIT[638*9 +: 8], INIT[637*9 +: 8], INIT[636*9 +: 8],
           INIT[635*9 +: 8], INIT[634*9 +: 8], INIT[633*9 +: 8], INIT[632*9 +: 8],
           INIT[631*9 +: 8], INIT[630*9 +: 8], INIT[629*9 +: 8], INIT[628*9 +: 8],
           INIT[627*9 +: 8], INIT[626*9 +: 8], INIT[625*9 +: 8], INIT[624*9 +: 8],
           INIT[623*9 +: 8], INIT[622*9 +: 8], INIT[621*9 +: 8], INIT[620*9 +: 8],
           INIT[619*9 +: 8], INIT[618*9 +: 8], INIT[617*9 +: 8], INIT[616*9 +: 8],
           INIT[615*9 +: 8], INIT[614*9 +: 8], INIT[613*9 +: 8], INIT[612*9 +: 8],
           INIT[611*9 +: 8], INIT[610*9 +: 8], INIT[609*9 +: 8], INIT[608*9 +: 8]}),
.INIT_14({ INIT[671*9 +: 8], INIT[670*9 +: 8], INIT[669*9 +: 8], INIT[668*9 +: 8],
           INIT[667*9 +: 8], INIT[666*9 +: 8], INIT[665*9 +: 8], INIT[664*9 +: 8],
           INIT[663*9 +: 8], INIT[662*9 +: 8], INIT[661*9 +: 8], INIT[660*9 +: 8],
           INIT[659*9 +: 8], INIT[658*9 +: 8], INIT[657*9 +: 8], INIT[656*9 +: 8],
           INIT[655*9 +: 8], INIT[654*9 +: 8], INIT[653*9 +: 8], INIT[652*9 +: 8],
           INIT[651*9 +: 8], INIT[650*9 +: 8], INIT[649*9 +: 8], INIT[648*9 +: 8],
           INIT[647*9 +: 8], INIT[646*9 +: 8], INIT[645*9 +: 8], INIT[644*9 +: 8],
           INIT[643*9 +: 8], INIT[642*9 +: 8], INIT[641*9 +: 8], INIT[640*9 +: 8]}),
.INIT_15({ INIT[703*9 +: 8], INIT[702*9 +: 8], INIT[701*9 +: 8], INIT[700*9 +: 8],
           INIT[699*9 +: 8], INIT[698*9 +: 8], INIT[697*9 +: 8], INIT[696*9 +: 8],
           INIT[695*9 +: 8], INIT[694*9 +: 8], INIT[693*9 +: 8], INIT[692*9 +: 8],
           INIT[691*9 +: 8], INIT[690*9 +: 8], INIT[689*9 +: 8], INIT[688*9 +: 8],
           INIT[687*9 +: 8], INIT[686*9 +: 8], INIT[685*9 +: 8], INIT[684*9 +: 8],
           INIT[683*9 +: 8], INIT[682*9 +: 8], INIT[681*9 +: 8], INIT[680*9 +: 8],
           INIT[679*9 +: 8], INIT[678*9 +: 8], INIT[677*9 +: 8], INIT[676*9 +: 8],
           INIT[675*9 +: 8], INIT[674*9 +: 8], INIT[673*9 +: 8], INIT[672*9 +: 8]}),
.INIT_16({ INIT[735*9 +: 8], INIT[734*9 +: 8], INIT[733*9 +: 8], INIT[732*9 +: 8],
           INIT[731*9 +: 8], INIT[730*9 +: 8], INIT[729*9 +: 8], INIT[728*9 +: 8],
           INIT[727*9 +: 8], INIT[726*9 +: 8], INIT[725*9 +: 8], INIT[724*9 +: 8],
           INIT[723*9 +: 8], INIT[722*9 +: 8], INIT[721*9 +: 8], INIT[720*9 +: 8],
           INIT[719*9 +: 8], INIT[718*9 +: 8], INIT[717*9 +: 8], INIT[716*9 +: 8],
           INIT[715*9 +: 8], INIT[714*9 +: 8], INIT[713*9 +: 8], INIT[712*9 +: 8],
           INIT[711*9 +: 8], INIT[710*9 +: 8], INIT[709*9 +: 8], INIT[708*9 +: 8],
           INIT[707*9 +: 8], INIT[706*9 +: 8], INIT[705*9 +: 8], INIT[704*9 +: 8]}),
.INIT_17({ INIT[767*9 +: 8], INIT[766*9 +: 8], INIT[765*9 +: 8], INIT[764*9 +: 8],
           INIT[763*9 +: 8], INIT[762*9 +: 8], INIT[761*9 +: 8], INIT[760*9 +: 8],
           INIT[759*9 +: 8], INIT[758*9 +: 8], INIT[757*9 +: 8], INIT[756*9 +: 8],
           INIT[755*9 +: 8], INIT[754*9 +: 8], INIT[753*9 +: 8], INIT[752*9 +: 8],
           INIT[751*9 +: 8], INIT[750*9 +: 8], INIT[749*9 +: 8], INIT[748*9 +: 8],
           INIT[747*9 +: 8], INIT[746*9 +: 8], INIT[745*9 +: 8], INIT[744*9 +: 8],
           INIT[743*9 +: 8], INIT[742*9 +: 8], INIT[741*9 +: 8], INIT[740*9 +: 8],
           INIT[739*9 +: 8], INIT[738*9 +: 8], INIT[737*9 +: 8], INIT[736*9 +: 8]}),
.INIT_18({ INIT[799*9 +: 8], INIT[798*9 +: 8], INIT[797*9 +: 8], INIT[796*9 +: 8],
           INIT[795*9 +: 8], INIT[794*9 +: 8], INIT[793*9 +: 8], INIT[792*9 +: 8],
           INIT[791*9 +: 8], INIT[790*9 +: 8], INIT[789*9 +: 8], INIT[788*9 +: 8],
           INIT[787*9 +: 8], INIT[786*9 +: 8], INIT[785*9 +: 8], INIT[784*9 +: 8],
           INIT[783*9 +: 8], INIT[782*9 +: 8], INIT[781*9 +: 8], INIT[780*9 +: 8],
           INIT[779*9 +: 8], INIT[778*9 +: 8], INIT[777*9 +: 8], INIT[776*9 +: 8],
           INIT[775*9 +: 8], INIT[774*9 +: 8], INIT[773*9 +: 8], INIT[772*9 +: 8],
           INIT[771*9 +: 8], INIT[770*9 +: 8], INIT[769*9 +: 8], INIT[768*9 +: 8]}),
.INIT_19({ INIT[831*9 +: 8], INIT[830*9 +: 8], INIT[829*9 +: 8], INIT[828*9 +: 8],
           INIT[827*9 +: 8], INIT[826*9 +: 8], INIT[825*9 +: 8], INIT[824*9 +: 8],
           INIT[823*9 +: 8], INIT[822*9 +: 8], INIT[821*9 +: 8], INIT[820*9 +: 8],
           INIT[819*9 +: 8], INIT[818*9 +: 8], INIT[817*9 +: 8], INIT[816*9 +: 8],
           INIT[815*9 +: 8], INIT[814*9 +: 8], INIT[813*9 +: 8], INIT[812*9 +: 8],
           INIT[811*9 +: 8], INIT[810*9 +: 8], INIT[809*9 +: 8], INIT[808*9 +: 8],
           INIT[807*9 +: 8], INIT[806*9 +: 8], INIT[805*9 +: 8], INIT[804*9 +: 8],
           INIT[803*9 +: 8], INIT[802*9 +: 8], INIT[801*9 +: 8], INIT[800*9 +: 8]}),
.INIT_1A({ INIT[863*9 +: 8], INIT[862*9 +: 8], INIT[861*9 +: 8], INIT[860*9 +: 8],
           INIT[859*9 +: 8], INIT[858*9 +: 8], INIT[857*9 +: 8], INIT[856*9 +: 8],
           INIT[855*9 +: 8], INIT[854*9 +: 8], INIT[853*9 +: 8], INIT[852*9 +: 8],
           INIT[851*9 +: 8], INIT[850*9 +: 8], INIT[849*9 +: 8], INIT[848*9 +: 8],
           INIT[847*9 +: 8], INIT[846*9 +: 8], INIT[845*9 +: 8], INIT[844*9 +: 8],
           INIT[843*9 +: 8], INIT[842*9 +: 8], INIT[841*9 +: 8], INIT[840*9 +: 8],
           INIT[839*9 +: 8], INIT[838*9 +: 8], INIT[837*9 +: 8], INIT[836*9 +: 8],
           INIT[835*9 +: 8], INIT[834*9 +: 8], INIT[833*9 +: 8], INIT[832*9 +: 8]}),
.INIT_1B({ INIT[895*9 +: 8], INIT[894*9 +: 8], INIT[893*9 +: 8], INIT[892*9 +: 8],
           INIT[891*9 +: 8], INIT[890*9 +: 8], INIT[889*9 +: 8], INIT[888*9 +: 8],
           INIT[887*9 +: 8], INIT[886*9 +: 8], INIT[885*9 +: 8], INIT[884*9 +: 8],
           INIT[883*9 +: 8], INIT[882*9 +: 8], INIT[881*9 +: 8], INIT[880*9 +: 8],
           INIT[879*9 +: 8], INIT[878*9 +: 8], INIT[877*9 +: 8], INIT[876*9 +: 8],
           INIT[875*9 +: 8], INIT[874*9 +: 8], INIT[873*9 +: 8], INIT[872*9 +: 8],
           INIT[871*9 +: 8], INIT[870*9 +: 8], INIT[869*9 +: 8], INIT[868*9 +: 8],
           INIT[867*9 +: 8], INIT[866*9 +: 8], INIT[865*9 +: 8], INIT[864*9 +: 8]}),
.INIT_1C({ INIT[927*9 +: 8], INIT[926*9 +: 8], INIT[925*9 +: 8], INIT[924*9 +: 8],
           INIT[923*9 +: 8], INIT[922*9 +: 8], INIT[921*9 +: 8], INIT[920*9 +: 8],
           INIT[919*9 +: 8], INIT[918*9 +: 8], INIT[917*9 +: 8], INIT[916*9 +: 8],
           INIT[915*9 +: 8], INIT[914*9 +: 8], INIT[913*9 +: 8], INIT[912*9 +: 8],
           INIT[911*9 +: 8], INIT[910*9 +: 8], INIT[909*9 +: 8], INIT[908*9 +: 8],
           INIT[907*9 +: 8], INIT[906*9 +: 8], INIT[905*9 +: 8], INIT[904*9 +: 8],
           INIT[903*9 +: 8], INIT[902*9 +: 8], INIT[901*9 +: 8], INIT[900*9 +: 8],
           INIT[899*9 +: 8], INIT[898*9 +: 8], INIT[897*9 +: 8], INIT[896*9 +: 8]}),
.INIT_1D({ INIT[959*9 +: 8], INIT[958*9 +: 8], INIT[957*9 +: 8], INIT[956*9 +: 8],
           INIT[955*9 +: 8], INIT[954*9 +: 8], INIT[953*9 +: 8], INIT[952*9 +: 8],
           INIT[951*9 +: 8], INIT[950*9 +: 8], INIT[949*9 +: 8], INIT[948*9 +: 8],
           INIT[947*9 +: 8], INIT[946*9 +: 8], INIT[945*9 +: 8], INIT[944*9 +: 8],
           INIT[943*9 +: 8], INIT[942*9 +: 8], INIT[941*9 +: 8], INIT[940*9 +: 8],
           INIT[939*9 +: 8], INIT[938*9 +: 8], INIT[937*9 +: 8], INIT[936*9 +: 8],
           INIT[935*9 +: 8], INIT[934*9 +: 8], INIT[933*9 +: 8], INIT[932*9 +: 8],
           INIT[931*9 +: 8], INIT[930*9 +: 8], INIT[929*9 +: 8], INIT[928*9 +: 8]}),
.INIT_1E({ INIT[991*9 +: 8], INIT[990*9 +: 8], INIT[989*9 +: 8], INIT[988*9 +: 8],
           INIT[987*9 +: 8], INIT[986*9 +: 8], INIT[985*9 +: 8], INIT[984*9 +: 8],
           INIT[983*9 +: 8], INIT[982*9 +: 8], INIT[981*9 +: 8], INIT[980*9 +: 8],
           INIT[979*9 +: 8], INIT[978*9 +: 8], INIT[977*9 +: 8], INIT[976*9 +: 8],
           INIT[975*9 +: 8], INIT[974*9 +: 8], INIT[973*9 +: 8], INIT[972*9 +: 8],
           INIT[971*9 +: 8], INIT[970*9 +: 8], INIT[969*9 +: 8], INIT[968*9 +: 8],
           INIT[967*9 +: 8], INIT[966*9 +: 8], INIT[965*9 +: 8], INIT[964*9 +: 8],
           INIT[963*9 +: 8], INIT[962*9 +: 8], INIT[961*9 +: 8], INIT[960*9 +: 8]}),
.INIT_1F({ INIT[1023*9 +: 8], INIT[1022*9 +: 8], INIT[1021*9 +: 8], INIT[1020*9 +: 8],
           INIT[1019*9 +: 8], INIT[1018*9 +: 8], INIT[1017*9 +: 8], INIT[1016*9 +: 8],
           INIT[1015*9 +: 8], INIT[1014*9 +: 8], INIT[1013*9 +: 8], INIT[1012*9 +: 8],
           INIT[1011*9 +: 8], INIT[1010*9 +: 8], INIT[1009*9 +: 8], INIT[1008*9 +: 8],
           INIT[1007*9 +: 8], INIT[1006*9 +: 8], INIT[1005*9 +: 8], INIT[1004*9 +: 8],
           INIT[1003*9 +: 8], INIT[1002*9 +: 8], INIT[1001*9 +: 8], INIT[1000*9 +: 8],
           INIT[999*9 +: 8], INIT[998*9 +: 8], INIT[997*9 +: 8], INIT[996*9 +: 8],
           INIT[995*9 +: 8], INIT[994*9 +: 8], INIT[993*9 +: 8], INIT[992*9 +: 8]}),
