    .ADA0(1'b0), .ADA1(1'b0), .ADA2(1'b0), .ADA3(A1ADDR[0]), .ADA4(A1ADDR[1]), .ADA5(A1ADDR[2]), .ADA6(A1ADDR[3]), .ADA7(A1ADDR[4]), .ADA8(A1ADDR[5]), .ADA9(A1ADDR[6]), .ADA10(A1ADDR[7]), .ADA11(A1ADDR[8]), .ADA12(A1ADDR[9]), .ADA13(A1ADDR[10]),
    .ADB0(1'b0), .ADB1(1'b0), .ADB2(1'b0), .ADB3(B1ADDR[0]), .ADB4(B1ADDR[1]), .ADB5(B1ADDR[2]), .ADB6(B1ADDR[3]), .ADB7(B1ADDR[4]), .ADB8(B1ADDR[5]), .ADB9(B1ADDR[6]), .ADB10(B1ADDR[7]), .ADB11(B1ADDR[8]), .ADB12(B1ADDR[9]), .ADB13(B1ADDR[10]),
    .DIA0(A1DATA[0]), .DIA1(A1DATA[1]), .DIA2(A1DATA[2]), .DIA3(A1DATA[3]), .DIA4(A1DATA[4]), .DIA5(A1DATA[5]), .DIA6(A1DATA[6]), .DIA7(A1DATA[7]), .DIA8(A1DATA[8]), .DIA9(1'b0), .DIA10(1'b0), .DIA11(1'b0), .DIA12(1'b0), .DIA13(1'b0), .DIA14(1'b0), .DIA15(1'b0), .DIA16(1'b0), .DIA17(1'b0),
    .DOB0(B1DATA[0]), .DOB1(B1DATA[1]), .DOB2(B1DATA[2]), .DOB3(B1DATA[3]), .DOB4(B1DATA[4]), .DOB5(B1DATA[5]), .DOB6(B1DATA[6]), .DOB7(B1DATA[7]), .DOB8(B1DATA[8]),
