    .ADA0(A1ADDR[0]), .ADA1(A1ADDR[1]), .ADA2(A1ADDR[2]), .ADA3(A1ADDR[3]), .ADA4(A1ADDR[4]), .ADA5(A1ADDR[5]), .ADA6(A1ADDR[6]), .ADA7(A1ADDR[7]), .ADA8(A1ADDR[8]), .ADA9(A1ADDR[9]), .ADA10(A1ADDR[10]), .ADA11(A1ADDR[11]), .ADA12(A1ADDR[12]), .ADA13(A1ADDR[13]),
    .ADB0(B1ADDR[0]), .ADB1(B1ADDR[1]), .ADB2(B1ADDR[2]), .ADB3(B1ADDR[3]), .ADB4(B1ADDR[4]), .ADB5(B1ADDR[5]), .ADB6(B1ADDR[6]), .ADB7(B1ADDR[7]), .ADB8(B1ADDR[8]), .ADB9(B1ADDR[9]), .ADB10(B1ADDR[10]), .ADB11(B1ADDR[11]), .ADB12(B1ADDR[12]), .ADB13(B1ADDR[13]),
    .DIA0(A1DATA[0]), .DIA1(1'b0), .DIA2(1'b0), .DIA3(1'b0), .DIA4(1'b0), .DIA5(1'b0), .DIA6(1'b0), .DIA7(1'b0), .DIA8(1'b0), .DIA9(1'b0), .DIA10(1'b0), .DIA11(1'b0), .DIA12(1'b0), .DIA13(1'b0), .DIA14(1'b0), .DIA15(1'b0), .DIA16(1'b0), .DIA17(1'b0),
    .DOB0(B1DATA[0]),
