    .ADW0(A1ADDR[0]), .ADW1(A1ADDR[1]), .ADW2(A1ADDR[2]), .ADW3(A1ADDR[3]), .ADW4(A1ADDR[4]), .ADW5(A1ADDR[5]), .ADW6(A1ADDR[6]), .ADW7(A1ADDR[7]), .ADW8(A1ADDR[8]),
    .ADR0(1'b0), .ADR1(1'b0), .ADR2(1'b0), .ADR3(1'b0), .ADR4(1'b0), .ADR5(B1ADDR[0]), .ADR6(B1ADDR[1]), .ADR7(B1ADDR[2]), .ADR8(B1ADDR[3]), .ADR9(B1ADDR[4]), .ADR10(B1ADDR[5]), .ADR11(B1ADDR[6]), .ADR12(B1ADDR[7]), .ADR13(B1ADDR[8]),
    .DI0(A1DATA[0]), .DI1(A1DATA[1]), .DI2(A1DATA[2]), .DI3(A1DATA[3]), .DI4(A1DATA[4]), .DI5(A1DATA[5]), .DI6(A1DATA[6]), .DI7(A1DATA[7]), .DI8(A1DATA[8]), .DI9(A1DATA[9]), .DI10(A1DATA[10]), .DI11(A1DATA[11]), .DI12(A1DATA[12]), .DI13(A1DATA[13]), .DI14(A1DATA[14]), .DI15(A1DATA[15]), .DI16(A1DATA[16]), .DI17(A1DATA[17]), .DI18(A1DATA[18]), .DI19(A1DATA[19]), .DI20(A1DATA[20]), .DI21(A1DATA[21]), .DI22(A1DATA[22]), .DI23(A1DATA[23]), .DI24(A1DATA[24]), .DI25(A1DATA[25]), .DI26(A1DATA[26]), .DI27(A1DATA[27]), .DI28(A1DATA[28]), .DI29(A1DATA[29]), .DI30(A1DATA[30]), .DI31(A1DATA[31]), .DI32(A1DATA[32]), .DI33(A1DATA[33]), .DI34(A1DATA[34]), .DI35(A1DATA[35]),
    .DO0(B1DATA[18]), .DO1(B1DATA[19]), .DO2(B1DATA[20]), .DO3(B1DATA[21]), .DO4(B1DATA[22]), .DO5(B1DATA[23]), .DO6(B1DATA[24]), .DO7(B1DATA[25]), .DO8(B1DATA[26]), .DO9(B1DATA[27]), .DO10(B1DATA[28]), .DO11(B1DATA[29]), .DO12(B1DATA[30]), .DO13(B1DATA[31]), .DO14(B1DATA[32]), .DO15(B1DATA[33]), .DO16(B1DATA[34]), .DO17(B1DATA[35]), .DO18(B1DATA[0]), .DO19(B1DATA[1]), .DO20(B1DATA[2]), .DO21(B1DATA[3]), .DO22(B1DATA[4]), .DO23(B1DATA[5]), .DO24(B1DATA[6]), .DO25(B1DATA[7]), .DO26(B1DATA[8]), .DO27(B1DATA[9]), .DO28(B1DATA[10]), .DO29(B1DATA[11]), .DO30(B1DATA[12]), .DO31(B1DATA[13]), .DO32(B1DATA[14]), .DO33(B1DATA[15]), .DO34(B1DATA[16]), .DO35(B1DATA[17]),
    .BE0(A1EN[0]), .BE1(A1EN[1]), .BE2(A1EN[2]), .BE3(A1EN[3]),
