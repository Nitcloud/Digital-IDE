.INITVAL_00({2'b00, INIT[ 15*18 +: 18], 2'b00, INIT[ 14*18 +: 18], 2'b00, INIT[ 13*18 +: 18], 2'b00, INIT[ 12*18 +: 18], 
          2'b00, INIT[ 11*18 +: 18], 2'b00, INIT[ 10*18 +: 18], 2'b00, INIT[  9*18 +: 18], 2'b00, INIT[  8*18 +: 18], 
          2'b00, INIT[  7*18 +: 18], 2'b00, INIT[  6*18 +: 18], 2'b00, INIT[  5*18 +: 18], 2'b00, INIT[  4*18 +: 18], 
          2'b00, INIT[  3*18 +: 18], 2'b00, INIT[  2*18 +: 18], 2'b00, INIT[  1*18 +: 18], 2'b00, INIT[  0*18 +: 18]}),
.INITVAL_01({2'b00, INIT[ 31*18 +: 18], 2'b00, INIT[ 30*18 +: 18], 2'b00, INIT[ 29*18 +: 18], 2'b00, INIT[ 28*18 +: 18], 
          2'b00, INIT[ 27*18 +: 18], 2'b00, INIT[ 26*18 +: 18], 2'b00, INIT[ 25*18 +: 18], 2'b00, INIT[ 24*18 +: 18], 
          2'b00, INIT[ 23*18 +: 18], 2'b00, INIT[ 22*18 +: 18], 2'b00, INIT[ 21*18 +: 18], 2'b00, INIT[ 20*18 +: 18], 
          2'b00, INIT[ 19*18 +: 18], 2'b00, INIT[ 18*18 +: 18], 2'b00, INIT[ 17*18 +: 18], 2'b00, INIT[ 16*18 +: 18]}),
.INITVAL_02({2'b00, INIT[ 47*18 +: 18], 2'b00, INIT[ 46*18 +: 18], 2'b00, INIT[ 45*18 +: 18], 2'b00, INIT[ 44*18 +: 18], 
          2'b00, INIT[ 43*18 +: 18], 2'b00, INIT[ 42*18 +: 18], 2'b00, INIT[ 41*18 +: 18], 2'b00, INIT[ 40*18 +: 18], 
          2'b00, INIT[ 39*18 +: 18], 2'b00, INIT[ 38*18 +: 18], 2'b00, INIT[ 37*18 +: 18], 2'b00, INIT[ 36*18 +: 18], 
          2'b00, INIT[ 35*18 +: 18], 2'b00, INIT[ 34*18 +: 18], 2'b00, INIT[ 33*18 +: 18], 2'b00, INIT[ 32*18 +: 18]}),
.INITVAL_03({2'b00, INIT[ 63*18 +: 18], 2'b00, INIT[ 62*18 +: 18], 2'b00, INIT[ 61*18 +: 18], 2'b00, INIT[ 60*18 +: 18], 
          2'b00, INIT[ 59*18 +: 18], 2'b00, INIT[ 58*18 +: 18], 2'b00, INIT[ 57*18 +: 18], 2'b00, INIT[ 56*18 +: 18], 
          2'b00, INIT[ 55*18 +: 18], 2'b00, INIT[ 54*18 +: 18], 2'b00, INIT[ 53*18 +: 18], 2'b00, INIT[ 52*18 +: 18], 
          2'b00, INIT[ 51*18 +: 18], 2'b00, INIT[ 50*18 +: 18], 2'b00, INIT[ 49*18 +: 18], 2'b00, INIT[ 48*18 +: 18]}),
.INITVAL_04({2'b00, INIT[ 79*18 +: 18], 2'b00, INIT[ 78*18 +: 18], 2'b00, INIT[ 77*18 +: 18], 2'b00, INIT[ 76*18 +: 18], 
          2'b00, INIT[ 75*18 +: 18], 2'b00, INIT[ 74*18 +: 18], 2'b00, INIT[ 73*18 +: 18], 2'b00, INIT[ 72*18 +: 18], 
          2'b00, INIT[ 71*18 +: 18], 2'b00, INIT[ 70*18 +: 18], 2'b00, INIT[ 69*18 +: 18], 2'b00, INIT[ 68*18 +: 18], 
          2'b00, INIT[ 67*18 +: 18], 2'b00, INIT[ 66*18 +: 18], 2'b00, INIT[ 65*18 +: 18], 2'b00, INIT[ 64*18 +: 18]}),
.INITVAL_05({2'b00, INIT[ 95*18 +: 18], 2'b00, INIT[ 94*18 +: 18], 2'b00, INIT[ 93*18 +: 18], 2'b00, INIT[ 92*18 +: 18], 
          2'b00, INIT[ 91*18 +: 18], 2'b00, INIT[ 90*18 +: 18], 2'b00, INIT[ 89*18 +: 18], 2'b00, INIT[ 88*18 +: 18], 
          2'b00, INIT[ 87*18 +: 18], 2'b00, INIT[ 86*18 +: 18], 2'b00, INIT[ 85*18 +: 18], 2'b00, INIT[ 84*18 +: 18], 
          2'b00, INIT[ 83*18 +: 18], 2'b00, INIT[ 82*18 +: 18], 2'b00, INIT[ 81*18 +: 18], 2'b00, INIT[ 80*18 +: 18]}),
.INITVAL_06({2'b00, INIT[111*18 +: 18], 2'b00, INIT[110*18 +: 18], 2'b00, INIT[109*18 +: 18], 2'b00, INIT[108*18 +: 18], 
          2'b00, INIT[107*18 +: 18], 2'b00, INIT[106*18 +: 18], 2'b00, INIT[105*18 +: 18], 2'b00, INIT[104*18 +: 18], 
          2'b00, INIT[103*18 +: 18], 2'b00, INIT[102*18 +: 18], 2'b00, INIT[101*18 +: 18], 2'b00, INIT[100*18 +: 18], 
          2'b00, INIT[ 99*18 +: 18], 2'b00, INIT[ 98*18 +: 18], 2'b00, INIT[ 97*18 +: 18], 2'b00, INIT[ 96*18 +: 18]}),
.INITVAL_07({2'b00, INIT[127*18 +: 18], 2'b00, INIT[126*18 +: 18], 2'b00, INIT[125*18 +: 18], 2'b00, INIT[124*18 +: 18], 
          2'b00, INIT[123*18 +: 18], 2'b00, INIT[122*18 +: 18], 2'b00, INIT[121*18 +: 18], 2'b00, INIT[120*18 +: 18], 
          2'b00, INIT[119*18 +: 18], 2'b00, INIT[118*18 +: 18], 2'b00, INIT[117*18 +: 18], 2'b00, INIT[116*18 +: 18], 
          2'b00, INIT[115*18 +: 18], 2'b00, INIT[114*18 +: 18], 2'b00, INIT[113*18 +: 18], 2'b00, INIT[112*18 +: 18]}),
.INITVAL_08({2'b00, INIT[143*18 +: 18], 2'b00, INIT[142*18 +: 18], 2'b00, INIT[141*18 +: 18], 2'b00, INIT[140*18 +: 18], 
          2'b00, INIT[139*18 +: 18], 2'b00, INIT[138*18 +: 18], 2'b00, INIT[137*18 +: 18], 2'b00, INIT[136*18 +: 18], 
          2'b00, INIT[135*18 +: 18], 2'b00, INIT[134*18 +: 18], 2'b00, INIT[133*18 +: 18], 2'b00, INIT[132*18 +: 18], 
          2'b00, INIT[131*18 +: 18], 2'b00, INIT[130*18 +: 18], 2'b00, INIT[129*18 +: 18], 2'b00, INIT[128*18 +: 18]}),
.INITVAL_09({2'b00, INIT[159*18 +: 18], 2'b00, INIT[158*18 +: 18], 2'b00, INIT[157*18 +: 18], 2'b00, INIT[156*18 +: 18], 
          2'b00, INIT[155*18 +: 18], 2'b00, INIT[154*18 +: 18], 2'b00, INIT[153*18 +: 18], 2'b00, INIT[152*18 +: 18], 
          2'b00, INIT[151*18 +: 18], 2'b00, INIT[150*18 +: 18], 2'b00, INIT[149*18 +: 18], 2'b00, INIT[148*18 +: 18], 
          2'b00, INIT[147*18 +: 18], 2'b00, INIT[146*18 +: 18], 2'b00, INIT[145*18 +: 18], 2'b00, INIT[144*18 +: 18]}),
.INITVAL_0A({2'b00, INIT[175*18 +: 18], 2'b00, INIT[174*18 +: 18], 2'b00, INIT[173*18 +: 18], 2'b00, INIT[172*18 +: 18], 
          2'b00, INIT[171*18 +: 18], 2'b00, INIT[170*18 +: 18], 2'b00, INIT[169*18 +: 18], 2'b00, INIT[168*18 +: 18], 
          2'b00, INIT[167*18 +: 18], 2'b00, INIT[166*18 +: 18], 2'b00, INIT[165*18 +: 18], 2'b00, INIT[164*18 +: 18], 
          2'b00, INIT[163*18 +: 18], 2'b00, INIT[162*18 +: 18], 2'b00, INIT[161*18 +: 18], 2'b00, INIT[160*18 +: 18]}),
.INITVAL_0B({2'b00, INIT[191*18 +: 18], 2'b00, INIT[190*18 +: 18], 2'b00, INIT[189*18 +: 18], 2'b00, INIT[188*18 +: 18], 
          2'b00, INIT[187*18 +: 18], 2'b00, INIT[186*18 +: 18], 2'b00, INIT[185*18 +: 18], 2'b00, INIT[184*18 +: 18], 
          2'b00, INIT[183*18 +: 18], 2'b00, INIT[182*18 +: 18], 2'b00, INIT[181*18 +: 18], 2'b00, INIT[180*18 +: 18], 
          2'b00, INIT[179*18 +: 18], 2'b00, INIT[178*18 +: 18], 2'b00, INIT[177*18 +: 18], 2'b00, INIT[176*18 +: 18]}),
.INITVAL_0C({2'b00, INIT[207*18 +: 18], 2'b00, INIT[206*18 +: 18], 2'b00, INIT[205*18 +: 18], 2'b00, INIT[204*18 +: 18], 
          2'b00, INIT[203*18 +: 18], 2'b00, INIT[202*18 +: 18], 2'b00, INIT[201*18 +: 18], 2'b00, INIT[200*18 +: 18], 
          2'b00, INIT[199*18 +: 18], 2'b00, INIT[198*18 +: 18], 2'b00, INIT[197*18 +: 18], 2'b00, INIT[196*18 +: 18], 
          2'b00, INIT[195*18 +: 18], 2'b00, INIT[194*18 +: 18], 2'b00, INIT[193*18 +: 18], 2'b00, INIT[192*18 +: 18]}),
.INITVAL_0D({2'b00, INIT[223*18 +: 18], 2'b00, INIT[222*18 +: 18], 2'b00, INIT[221*18 +: 18], 2'b00, INIT[220*18 +: 18], 
          2'b00, INIT[219*18 +: 18], 2'b00, INIT[218*18 +: 18], 2'b00, INIT[217*18 +: 18], 2'b00, INIT[216*18 +: 18], 
          2'b00, INIT[215*18 +: 18], 2'b00, INIT[214*18 +: 18], 2'b00, INIT[213*18 +: 18], 2'b00, INIT[212*18 +: 18], 
          2'b00, INIT[211*18 +: 18], 2'b00, INIT[210*18 +: 18], 2'b00, INIT[209*18 +: 18], 2'b00, INIT[208*18 +: 18]}),
.INITVAL_0E({2'b00, INIT[239*18 +: 18], 2'b00, INIT[238*18 +: 18], 2'b00, INIT[237*18 +: 18], 2'b00, INIT[236*18 +: 18], 
          2'b00, INIT[235*18 +: 18], 2'b00, INIT[234*18 +: 18], 2'b00, INIT[233*18 +: 18], 2'b00, INIT[232*18 +: 18], 
          2'b00, INIT[231*18 +: 18], 2'b00, INIT[230*18 +: 18], 2'b00, INIT[229*18 +: 18], 2'b00, INIT[228*18 +: 18], 
          2'b00, INIT[227*18 +: 18], 2'b00, INIT[226*18 +: 18], 2'b00, INIT[225*18 +: 18], 2'b00, INIT[224*18 +: 18]}),
.INITVAL_0F({2'b00, INIT[255*18 +: 18], 2'b00, INIT[254*18 +: 18], 2'b00, INIT[253*18 +: 18], 2'b00, INIT[252*18 +: 18], 
          2'b00, INIT[251*18 +: 18], 2'b00, INIT[250*18 +: 18], 2'b00, INIT[249*18 +: 18], 2'b00, INIT[248*18 +: 18], 
          2'b00, INIT[247*18 +: 18], 2'b00, INIT[246*18 +: 18], 2'b00, INIT[245*18 +: 18], 2'b00, INIT[244*18 +: 18], 
          2'b00, INIT[243*18 +: 18], 2'b00, INIT[242*18 +: 18], 2'b00, INIT[241*18 +: 18], 2'b00, INIT[240*18 +: 18]}),
.INITVAL_10({2'b00, INIT[271*18 +: 18], 2'b00, INIT[270*18 +: 18], 2'b00, INIT[269*18 +: 18], 2'b00, INIT[268*18 +: 18], 
          2'b00, INIT[267*18 +: 18], 2'b00, INIT[266*18 +: 18], 2'b00, INIT[265*18 +: 18], 2'b00, INIT[264*18 +: 18], 
          2'b00, INIT[263*18 +: 18], 2'b00, INIT[262*18 +: 18], 2'b00, INIT[261*18 +: 18], 2'b00, INIT[260*18 +: 18], 
          2'b00, INIT[259*18 +: 18], 2'b00, INIT[258*18 +: 18], 2'b00, INIT[257*18 +: 18], 2'b00, INIT[256*18 +: 18]}),
.INITVAL_11({2'b00, INIT[287*18 +: 18], 2'b00, INIT[286*18 +: 18], 2'b00, INIT[285*18 +: 18], 2'b00, INIT[284*18 +: 18], 
          2'b00, INIT[283*18 +: 18], 2'b00, INIT[282*18 +: 18], 2'b00, INIT[281*18 +: 18], 2'b00, INIT[280*18 +: 18], 
          2'b00, INIT[279*18 +: 18], 2'b00, INIT[278*18 +: 18], 2'b00, INIT[277*18 +: 18], 2'b00, INIT[276*18 +: 18], 
          2'b00, INIT[275*18 +: 18], 2'b00, INIT[274*18 +: 18], 2'b00, INIT[273*18 +: 18], 2'b00, INIT[272*18 +: 18]}),
.INITVAL_12({2'b00, INIT[303*18 +: 18], 2'b00, INIT[302*18 +: 18], 2'b00, INIT[301*18 +: 18], 2'b00, INIT[300*18 +: 18], 
          2'b00, INIT[299*18 +: 18], 2'b00, INIT[298*18 +: 18], 2'b00, INIT[297*18 +: 18], 2'b00, INIT[296*18 +: 18], 
          2'b00, INIT[295*18 +: 18], 2'b00, INIT[294*18 +: 18], 2'b00, INIT[293*18 +: 18], 2'b00, INIT[292*18 +: 18], 
          2'b00, INIT[291*18 +: 18], 2'b00, INIT[290*18 +: 18], 2'b00, INIT[289*18 +: 18], 2'b00, INIT[288*18 +: 18]}),
.INITVAL_13({2'b00, INIT[319*18 +: 18], 2'b00, INIT[318*18 +: 18], 2'b00, INIT[317*18 +: 18], 2'b00, INIT[316*18 +: 18], 
          2'b00, INIT[315*18 +: 18], 2'b00, INIT[314*18 +: 18], 2'b00, INIT[313*18 +: 18], 2'b00, INIT[312*18 +: 18], 
          2'b00, INIT[311*18 +: 18], 2'b00, INIT[310*18 +: 18], 2'b00, INIT[309*18 +: 18], 2'b00, INIT[308*18 +: 18], 
          2'b00, INIT[307*18 +: 18], 2'b00, INIT[306*18 +: 18], 2'b00, INIT[305*18 +: 18], 2'b00, INIT[304*18 +: 18]}),
.INITVAL_14({2'b00, INIT[335*18 +: 18], 2'b00, INIT[334*18 +: 18], 2'b00, INIT[333*18 +: 18], 2'b00, INIT[332*18 +: 18], 
          2'b00, INIT[331*18 +: 18], 2'b00, INIT[330*18 +: 18], 2'b00, INIT[329*18 +: 18], 2'b00, INIT[328*18 +: 18], 
          2'b00, INIT[327*18 +: 18], 2'b00, INIT[326*18 +: 18], 2'b00, INIT[325*18 +: 18], 2'b00, INIT[324*18 +: 18], 
          2'b00, INIT[323*18 +: 18], 2'b00, INIT[322*18 +: 18], 2'b00, INIT[321*18 +: 18], 2'b00, INIT[320*18 +: 18]}),
.INITVAL_15({2'b00, INIT[351*18 +: 18], 2'b00, INIT[350*18 +: 18], 2'b00, INIT[349*18 +: 18], 2'b00, INIT[348*18 +: 18], 
          2'b00, INIT[347*18 +: 18], 2'b00, INIT[346*18 +: 18], 2'b00, INIT[345*18 +: 18], 2'b00, INIT[344*18 +: 18], 
          2'b00, INIT[343*18 +: 18], 2'b00, INIT[342*18 +: 18], 2'b00, INIT[341*18 +: 18], 2'b00, INIT[340*18 +: 18], 
          2'b00, INIT[339*18 +: 18], 2'b00, INIT[338*18 +: 18], 2'b00, INIT[337*18 +: 18], 2'b00, INIT[336*18 +: 18]}),
.INITVAL_16({2'b00, INIT[367*18 +: 18], 2'b00, INIT[366*18 +: 18], 2'b00, INIT[365*18 +: 18], 2'b00, INIT[364*18 +: 18], 
          2'b00, INIT[363*18 +: 18], 2'b00, INIT[362*18 +: 18], 2'b00, INIT[361*18 +: 18], 2'b00, INIT[360*18 +: 18], 
          2'b00, INIT[359*18 +: 18], 2'b00, INIT[358*18 +: 18], 2'b00, INIT[357*18 +: 18], 2'b00, INIT[356*18 +: 18], 
          2'b00, INIT[355*18 +: 18], 2'b00, INIT[354*18 +: 18], 2'b00, INIT[353*18 +: 18], 2'b00, INIT[352*18 +: 18]}),
.INITVAL_17({2'b00, INIT[383*18 +: 18], 2'b00, INIT[382*18 +: 18], 2'b00, INIT[381*18 +: 18], 2'b00, INIT[380*18 +: 18], 
          2'b00, INIT[379*18 +: 18], 2'b00, INIT[378*18 +: 18], 2'b00, INIT[377*18 +: 18], 2'b00, INIT[376*18 +: 18], 
          2'b00, INIT[375*18 +: 18], 2'b00, INIT[374*18 +: 18], 2'b00, INIT[373*18 +: 18], 2'b00, INIT[372*18 +: 18], 
          2'b00, INIT[371*18 +: 18], 2'b00, INIT[370*18 +: 18], 2'b00, INIT[369*18 +: 18], 2'b00, INIT[368*18 +: 18]}),
.INITVAL_18({2'b00, INIT[399*18 +: 18], 2'b00, INIT[398*18 +: 18], 2'b00, INIT[397*18 +: 18], 2'b00, INIT[396*18 +: 18], 
          2'b00, INIT[395*18 +: 18], 2'b00, INIT[394*18 +: 18], 2'b00, INIT[393*18 +: 18], 2'b00, INIT[392*18 +: 18], 
          2'b00, INIT[391*18 +: 18], 2'b00, INIT[390*18 +: 18], 2'b00, INIT[389*18 +: 18], 2'b00, INIT[388*18 +: 18], 
          2'b00, INIT[387*18 +: 18], 2'b00, INIT[386*18 +: 18], 2'b00, INIT[385*18 +: 18], 2'b00, INIT[384*18 +: 18]}),
.INITVAL_19({2'b00, INIT[415*18 +: 18], 2'b00, INIT[414*18 +: 18], 2'b00, INIT[413*18 +: 18], 2'b00, INIT[412*18 +: 18], 
          2'b00, INIT[411*18 +: 18], 2'b00, INIT[410*18 +: 18], 2'b00, INIT[409*18 +: 18], 2'b00, INIT[408*18 +: 18], 
          2'b00, INIT[407*18 +: 18], 2'b00, INIT[406*18 +: 18], 2'b00, INIT[405*18 +: 18], 2'b00, INIT[404*18 +: 18], 
          2'b00, INIT[403*18 +: 18], 2'b00, INIT[402*18 +: 18], 2'b00, INIT[401*18 +: 18], 2'b00, INIT[400*18 +: 18]}),
.INITVAL_1A({2'b00, INIT[431*18 +: 18], 2'b00, INIT[430*18 +: 18], 2'b00, INIT[429*18 +: 18], 2'b00, INIT[428*18 +: 18], 
          2'b00, INIT[427*18 +: 18], 2'b00, INIT[426*18 +: 18], 2'b00, INIT[425*18 +: 18], 2'b00, INIT[424*18 +: 18], 
          2'b00, INIT[423*18 +: 18], 2'b00, INIT[422*18 +: 18], 2'b00, INIT[421*18 +: 18], 2'b00, INIT[420*18 +: 18], 
          2'b00, INIT[419*18 +: 18], 2'b00, INIT[418*18 +: 18], 2'b00, INIT[417*18 +: 18], 2'b00, INIT[416*18 +: 18]}),
.INITVAL_1B({2'b00, INIT[447*18 +: 18], 2'b00, INIT[446*18 +: 18], 2'b00, INIT[445*18 +: 18], 2'b00, INIT[444*18 +: 18], 
          2'b00, INIT[443*18 +: 18], 2'b00, INIT[442*18 +: 18], 2'b00, INIT[441*18 +: 18], 2'b00, INIT[440*18 +: 18], 
          2'b00, INIT[439*18 +: 18], 2'b00, INIT[438*18 +: 18], 2'b00, INIT[437*18 +: 18], 2'b00, INIT[436*18 +: 18], 
          2'b00, INIT[435*18 +: 18], 2'b00, INIT[434*18 +: 18], 2'b00, INIT[433*18 +: 18], 2'b00, INIT[432*18 +: 18]}),
.INITVAL_1C({2'b00, INIT[463*18 +: 18], 2'b00, INIT[462*18 +: 18], 2'b00, INIT[461*18 +: 18], 2'b00, INIT[460*18 +: 18], 
          2'b00, INIT[459*18 +: 18], 2'b00, INIT[458*18 +: 18], 2'b00, INIT[457*18 +: 18], 2'b00, INIT[456*18 +: 18], 
          2'b00, INIT[455*18 +: 18], 2'b00, INIT[454*18 +: 18], 2'b00, INIT[453*18 +: 18], 2'b00, INIT[452*18 +: 18], 
          2'b00, INIT[451*18 +: 18], 2'b00, INIT[450*18 +: 18], 2'b00, INIT[449*18 +: 18], 2'b00, INIT[448*18 +: 18]}),
.INITVAL_1D({2'b00, INIT[479*18 +: 18], 2'b00, INIT[478*18 +: 18], 2'b00, INIT[477*18 +: 18], 2'b00, INIT[476*18 +: 18], 
          2'b00, INIT[475*18 +: 18], 2'b00, INIT[474*18 +: 18], 2'b00, INIT[473*18 +: 18], 2'b00, INIT[472*18 +: 18], 
          2'b00, INIT[471*18 +: 18], 2'b00, INIT[470*18 +: 18], 2'b00, INIT[469*18 +: 18], 2'b00, INIT[468*18 +: 18], 
          2'b00, INIT[467*18 +: 18], 2'b00, INIT[466*18 +: 18], 2'b00, INIT[465*18 +: 18], 2'b00, INIT[464*18 +: 18]}),
.INITVAL_1E({2'b00, INIT[495*18 +: 18], 2'b00, INIT[494*18 +: 18], 2'b00, INIT[493*18 +: 18], 2'b00, INIT[492*18 +: 18], 
          2'b00, INIT[491*18 +: 18], 2'b00, INIT[490*18 +: 18], 2'b00, INIT[489*18 +: 18], 2'b00, INIT[488*18 +: 18], 
          2'b00, INIT[487*18 +: 18], 2'b00, INIT[486*18 +: 18], 2'b00, INIT[485*18 +: 18], 2'b00, INIT[484*18 +: 18], 
          2'b00, INIT[483*18 +: 18], 2'b00, INIT[482*18 +: 18], 2'b00, INIT[481*18 +: 18], 2'b00, INIT[480*18 +: 18]}),
.INITVAL_1F({2'b00, INIT[511*18 +: 18], 2'b00, INIT[510*18 +: 18], 2'b00, INIT[509*18 +: 18], 2'b00, INIT[508*18 +: 18], 
          2'b00, INIT[507*18 +: 18], 2'b00, INIT[506*18 +: 18], 2'b00, INIT[505*18 +: 18], 2'b00, INIT[504*18 +: 18], 
          2'b00, INIT[503*18 +: 18], 2'b00, INIT[502*18 +: 18], 2'b00, INIT[501*18 +: 18], 2'b00, INIT[500*18 +: 18], 
          2'b00, INIT[499*18 +: 18], 2'b00, INIT[498*18 +: 18], 2'b00, INIT[497*18 +: 18], 2'b00, INIT[496*18 +: 18]}),
.INITVAL_20({2'b00, INIT[527*18 +: 18], 2'b00, INIT[526*18 +: 18], 2'b00, INIT[525*18 +: 18], 2'b00, INIT[524*18 +: 18], 
          2'b00, INIT[523*18 +: 18], 2'b00, INIT[522*18 +: 18], 2'b00, INIT[521*18 +: 18], 2'b00, INIT[520*18 +: 18], 
          2'b00, INIT[519*18 +: 18], 2'b00, INIT[518*18 +: 18], 2'b00, INIT[517*18 +: 18], 2'b00, INIT[516*18 +: 18], 
          2'b00, INIT[515*18 +: 18], 2'b00, INIT[514*18 +: 18], 2'b00, INIT[513*18 +: 18], 2'b00, INIT[512*18 +: 18]}),
.INITVAL_21({2'b00, INIT[543*18 +: 18], 2'b00, INIT[542*18 +: 18], 2'b00, INIT[541*18 +: 18], 2'b00, INIT[540*18 +: 18], 
          2'b00, INIT[539*18 +: 18], 2'b00, INIT[538*18 +: 18], 2'b00, INIT[537*18 +: 18], 2'b00, INIT[536*18 +: 18], 
          2'b00, INIT[535*18 +: 18], 2'b00, INIT[534*18 +: 18], 2'b00, INIT[533*18 +: 18], 2'b00, INIT[532*18 +: 18], 
          2'b00, INIT[531*18 +: 18], 2'b00, INIT[530*18 +: 18], 2'b00, INIT[529*18 +: 18], 2'b00, INIT[528*18 +: 18]}),
.INITVAL_22({2'b00, INIT[559*18 +: 18], 2'b00, INIT[558*18 +: 18], 2'b00, INIT[557*18 +: 18], 2'b00, INIT[556*18 +: 18], 
          2'b00, INIT[555*18 +: 18], 2'b00, INIT[554*18 +: 18], 2'b00, INIT[553*18 +: 18], 2'b00, INIT[552*18 +: 18], 
          2'b00, INIT[551*18 +: 18], 2'b00, INIT[550*18 +: 18], 2'b00, INIT[549*18 +: 18], 2'b00, INIT[548*18 +: 18], 
          2'b00, INIT[547*18 +: 18], 2'b00, INIT[546*18 +: 18], 2'b00, INIT[545*18 +: 18], 2'b00, INIT[544*18 +: 18]}),
.INITVAL_23({2'b00, INIT[575*18 +: 18], 2'b00, INIT[574*18 +: 18], 2'b00, INIT[573*18 +: 18], 2'b00, INIT[572*18 +: 18], 
          2'b00, INIT[571*18 +: 18], 2'b00, INIT[570*18 +: 18], 2'b00, INIT[569*18 +: 18], 2'b00, INIT[568*18 +: 18], 
          2'b00, INIT[567*18 +: 18], 2'b00, INIT[566*18 +: 18], 2'b00, INIT[565*18 +: 18], 2'b00, INIT[564*18 +: 18], 
          2'b00, INIT[563*18 +: 18], 2'b00, INIT[562*18 +: 18], 2'b00, INIT[561*18 +: 18], 2'b00, INIT[560*18 +: 18]}),
.INITVAL_24({2'b00, INIT[591*18 +: 18], 2'b00, INIT[590*18 +: 18], 2'b00, INIT[589*18 +: 18], 2'b00, INIT[588*18 +: 18], 
          2'b00, INIT[587*18 +: 18], 2'b00, INIT[586*18 +: 18], 2'b00, INIT[585*18 +: 18], 2'b00, INIT[584*18 +: 18], 
          2'b00, INIT[583*18 +: 18], 2'b00, INIT[582*18 +: 18], 2'b00, INIT[581*18 +: 18], 2'b00, INIT[580*18 +: 18], 
          2'b00, INIT[579*18 +: 18], 2'b00, INIT[578*18 +: 18], 2'b00, INIT[577*18 +: 18], 2'b00, INIT[576*18 +: 18]}),
.INITVAL_25({2'b00, INIT[607*18 +: 18], 2'b00, INIT[606*18 +: 18], 2'b00, INIT[605*18 +: 18], 2'b00, INIT[604*18 +: 18], 
          2'b00, INIT[603*18 +: 18], 2'b00, INIT[602*18 +: 18], 2'b00, INIT[601*18 +: 18], 2'b00, INIT[600*18 +: 18], 
          2'b00, INIT[599*18 +: 18], 2'b00, INIT[598*18 +: 18], 2'b00, INIT[597*18 +: 18], 2'b00, INIT[596*18 +: 18], 
          2'b00, INIT[595*18 +: 18], 2'b00, INIT[594*18 +: 18], 2'b00, INIT[593*18 +: 18], 2'b00, INIT[592*18 +: 18]}),
.INITVAL_26({2'b00, INIT[623*18 +: 18], 2'b00, INIT[622*18 +: 18], 2'b00, INIT[621*18 +: 18], 2'b00, INIT[620*18 +: 18], 
          2'b00, INIT[619*18 +: 18], 2'b00, INIT[618*18 +: 18], 2'b00, INIT[617*18 +: 18], 2'b00, INIT[616*18 +: 18], 
          2'b00, INIT[615*18 +: 18], 2'b00, INIT[614*18 +: 18], 2'b00, INIT[613*18 +: 18], 2'b00, INIT[612*18 +: 18], 
          2'b00, INIT[611*18 +: 18], 2'b00, INIT[610*18 +: 18], 2'b00, INIT[609*18 +: 18], 2'b00, INIT[608*18 +: 18]}),
.INITVAL_27({2'b00, INIT[639*18 +: 18], 2'b00, INIT[638*18 +: 18], 2'b00, INIT[637*18 +: 18], 2'b00, INIT[636*18 +: 18], 
          2'b00, INIT[635*18 +: 18], 2'b00, INIT[634*18 +: 18], 2'b00, INIT[633*18 +: 18], 2'b00, INIT[632*18 +: 18], 
          2'b00, INIT[631*18 +: 18], 2'b00, INIT[630*18 +: 18], 2'b00, INIT[629*18 +: 18], 2'b00, INIT[628*18 +: 18], 
          2'b00, INIT[627*18 +: 18], 2'b00, INIT[626*18 +: 18], 2'b00, INIT[625*18 +: 18], 2'b00, INIT[624*18 +: 18]}),
.INITVAL_28({2'b00, INIT[655*18 +: 18], 2'b00, INIT[654*18 +: 18], 2'b00, INIT[653*18 +: 18], 2'b00, INIT[652*18 +: 18], 
          2'b00, INIT[651*18 +: 18], 2'b00, INIT[650*18 +: 18], 2'b00, INIT[649*18 +: 18], 2'b00, INIT[648*18 +: 18], 
          2'b00, INIT[647*18 +: 18], 2'b00, INIT[646*18 +: 18], 2'b00, INIT[645*18 +: 18], 2'b00, INIT[644*18 +: 18], 
          2'b00, INIT[643*18 +: 18], 2'b00, INIT[642*18 +: 18], 2'b00, INIT[641*18 +: 18], 2'b00, INIT[640*18 +: 18]}),
.INITVAL_29({2'b00, INIT[671*18 +: 18], 2'b00, INIT[670*18 +: 18], 2'b00, INIT[669*18 +: 18], 2'b00, INIT[668*18 +: 18], 
          2'b00, INIT[667*18 +: 18], 2'b00, INIT[666*18 +: 18], 2'b00, INIT[665*18 +: 18], 2'b00, INIT[664*18 +: 18], 
          2'b00, INIT[663*18 +: 18], 2'b00, INIT[662*18 +: 18], 2'b00, INIT[661*18 +: 18], 2'b00, INIT[660*18 +: 18], 
          2'b00, INIT[659*18 +: 18], 2'b00, INIT[658*18 +: 18], 2'b00, INIT[657*18 +: 18], 2'b00, INIT[656*18 +: 18]}),
.INITVAL_2A({2'b00, INIT[687*18 +: 18], 2'b00, INIT[686*18 +: 18], 2'b00, INIT[685*18 +: 18], 2'b00, INIT[684*18 +: 18], 
          2'b00, INIT[683*18 +: 18], 2'b00, INIT[682*18 +: 18], 2'b00, INIT[681*18 +: 18], 2'b00, INIT[680*18 +: 18], 
          2'b00, INIT[679*18 +: 18], 2'b00, INIT[678*18 +: 18], 2'b00, INIT[677*18 +: 18], 2'b00, INIT[676*18 +: 18], 
          2'b00, INIT[675*18 +: 18], 2'b00, INIT[674*18 +: 18], 2'b00, INIT[673*18 +: 18], 2'b00, INIT[672*18 +: 18]}),
.INITVAL_2B({2'b00, INIT[703*18 +: 18], 2'b00, INIT[702*18 +: 18], 2'b00, INIT[701*18 +: 18], 2'b00, INIT[700*18 +: 18], 
          2'b00, INIT[699*18 +: 18], 2'b00, INIT[698*18 +: 18], 2'b00, INIT[697*18 +: 18], 2'b00, INIT[696*18 +: 18], 
          2'b00, INIT[695*18 +: 18], 2'b00, INIT[694*18 +: 18], 2'b00, INIT[693*18 +: 18], 2'b00, INIT[692*18 +: 18], 
          2'b00, INIT[691*18 +: 18], 2'b00, INIT[690*18 +: 18], 2'b00, INIT[689*18 +: 18], 2'b00, INIT[688*18 +: 18]}),
.INITVAL_2C({2'b00, INIT[719*18 +: 18], 2'b00, INIT[718*18 +: 18], 2'b00, INIT[717*18 +: 18], 2'b00, INIT[716*18 +: 18], 
          2'b00, INIT[715*18 +: 18], 2'b00, INIT[714*18 +: 18], 2'b00, INIT[713*18 +: 18], 2'b00, INIT[712*18 +: 18], 
          2'b00, INIT[711*18 +: 18], 2'b00, INIT[710*18 +: 18], 2'b00, INIT[709*18 +: 18], 2'b00, INIT[708*18 +: 18], 
          2'b00, INIT[707*18 +: 18], 2'b00, INIT[706*18 +: 18], 2'b00, INIT[705*18 +: 18], 2'b00, INIT[704*18 +: 18]}),
.INITVAL_2D({2'b00, INIT[735*18 +: 18], 2'b00, INIT[734*18 +: 18], 2'b00, INIT[733*18 +: 18], 2'b00, INIT[732*18 +: 18], 
          2'b00, INIT[731*18 +: 18], 2'b00, INIT[730*18 +: 18], 2'b00, INIT[729*18 +: 18], 2'b00, INIT[728*18 +: 18], 
          2'b00, INIT[727*18 +: 18], 2'b00, INIT[726*18 +: 18], 2'b00, INIT[725*18 +: 18], 2'b00, INIT[724*18 +: 18], 
          2'b00, INIT[723*18 +: 18], 2'b00, INIT[722*18 +: 18], 2'b00, INIT[721*18 +: 18], 2'b00, INIT[720*18 +: 18]}),
.INITVAL_2E({2'b00, INIT[751*18 +: 18], 2'b00, INIT[750*18 +: 18], 2'b00, INIT[749*18 +: 18], 2'b00, INIT[748*18 +: 18], 
          2'b00, INIT[747*18 +: 18], 2'b00, INIT[746*18 +: 18], 2'b00, INIT[745*18 +: 18], 2'b00, INIT[744*18 +: 18], 
          2'b00, INIT[743*18 +: 18], 2'b00, INIT[742*18 +: 18], 2'b00, INIT[741*18 +: 18], 2'b00, INIT[740*18 +: 18], 
          2'b00, INIT[739*18 +: 18], 2'b00, INIT[738*18 +: 18], 2'b00, INIT[737*18 +: 18], 2'b00, INIT[736*18 +: 18]}),
.INITVAL_2F({2'b00, INIT[767*18 +: 18], 2'b00, INIT[766*18 +: 18], 2'b00, INIT[765*18 +: 18], 2'b00, INIT[764*18 +: 18], 
          2'b00, INIT[763*18 +: 18], 2'b00, INIT[762*18 +: 18], 2'b00, INIT[761*18 +: 18], 2'b00, INIT[760*18 +: 18], 
          2'b00, INIT[759*18 +: 18], 2'b00, INIT[758*18 +: 18], 2'b00, INIT[757*18 +: 18], 2'b00, INIT[756*18 +: 18], 
          2'b00, INIT[755*18 +: 18], 2'b00, INIT[754*18 +: 18], 2'b00, INIT[753*18 +: 18], 2'b00, INIT[752*18 +: 18]}),
.INITVAL_30({2'b00, INIT[783*18 +: 18], 2'b00, INIT[782*18 +: 18], 2'b00, INIT[781*18 +: 18], 2'b00, INIT[780*18 +: 18], 
          2'b00, INIT[779*18 +: 18], 2'b00, INIT[778*18 +: 18], 2'b00, INIT[777*18 +: 18], 2'b00, INIT[776*18 +: 18], 
          2'b00, INIT[775*18 +: 18], 2'b00, INIT[774*18 +: 18], 2'b00, INIT[773*18 +: 18], 2'b00, INIT[772*18 +: 18], 
          2'b00, INIT[771*18 +: 18], 2'b00, INIT[770*18 +: 18], 2'b00, INIT[769*18 +: 18], 2'b00, INIT[768*18 +: 18]}),
.INITVAL_31({2'b00, INIT[799*18 +: 18], 2'b00, INIT[798*18 +: 18], 2'b00, INIT[797*18 +: 18], 2'b00, INIT[796*18 +: 18], 
          2'b00, INIT[795*18 +: 18], 2'b00, INIT[794*18 +: 18], 2'b00, INIT[793*18 +: 18], 2'b00, INIT[792*18 +: 18], 
          2'b00, INIT[791*18 +: 18], 2'b00, INIT[790*18 +: 18], 2'b00, INIT[789*18 +: 18], 2'b00, INIT[788*18 +: 18], 
          2'b00, INIT[787*18 +: 18], 2'b00, INIT[786*18 +: 18], 2'b00, INIT[785*18 +: 18], 2'b00, INIT[784*18 +: 18]}),
.INITVAL_32({2'b00, INIT[815*18 +: 18], 2'b00, INIT[814*18 +: 18], 2'b00, INIT[813*18 +: 18], 2'b00, INIT[812*18 +: 18], 
          2'b00, INIT[811*18 +: 18], 2'b00, INIT[810*18 +: 18], 2'b00, INIT[809*18 +: 18], 2'b00, INIT[808*18 +: 18], 
          2'b00, INIT[807*18 +: 18], 2'b00, INIT[806*18 +: 18], 2'b00, INIT[805*18 +: 18], 2'b00, INIT[804*18 +: 18], 
          2'b00, INIT[803*18 +: 18], 2'b00, INIT[802*18 +: 18], 2'b00, INIT[801*18 +: 18], 2'b00, INIT[800*18 +: 18]}),
.INITVAL_33({2'b00, INIT[831*18 +: 18], 2'b00, INIT[830*18 +: 18], 2'b00, INIT[829*18 +: 18], 2'b00, INIT[828*18 +: 18], 
          2'b00, INIT[827*18 +: 18], 2'b00, INIT[826*18 +: 18], 2'b00, INIT[825*18 +: 18], 2'b00, INIT[824*18 +: 18], 
          2'b00, INIT[823*18 +: 18], 2'b00, INIT[822*18 +: 18], 2'b00, INIT[821*18 +: 18], 2'b00, INIT[820*18 +: 18], 
          2'b00, INIT[819*18 +: 18], 2'b00, INIT[818*18 +: 18], 2'b00, INIT[817*18 +: 18], 2'b00, INIT[816*18 +: 18]}),
.INITVAL_34({2'b00, INIT[847*18 +: 18], 2'b00, INIT[846*18 +: 18], 2'b00, INIT[845*18 +: 18], 2'b00, INIT[844*18 +: 18], 
          2'b00, INIT[843*18 +: 18], 2'b00, INIT[842*18 +: 18], 2'b00, INIT[841*18 +: 18], 2'b00, INIT[840*18 +: 18], 
          2'b00, INIT[839*18 +: 18], 2'b00, INIT[838*18 +: 18], 2'b00, INIT[837*18 +: 18], 2'b00, INIT[836*18 +: 18], 
          2'b00, INIT[835*18 +: 18], 2'b00, INIT[834*18 +: 18], 2'b00, INIT[833*18 +: 18], 2'b00, INIT[832*18 +: 18]}),
.INITVAL_35({2'b00, INIT[863*18 +: 18], 2'b00, INIT[862*18 +: 18], 2'b00, INIT[861*18 +: 18], 2'b00, INIT[860*18 +: 18], 
          2'b00, INIT[859*18 +: 18], 2'b00, INIT[858*18 +: 18], 2'b00, INIT[857*18 +: 18], 2'b00, INIT[856*18 +: 18], 
          2'b00, INIT[855*18 +: 18], 2'b00, INIT[854*18 +: 18], 2'b00, INIT[853*18 +: 18], 2'b00, INIT[852*18 +: 18], 
          2'b00, INIT[851*18 +: 18], 2'b00, INIT[850*18 +: 18], 2'b00, INIT[849*18 +: 18], 2'b00, INIT[848*18 +: 18]}),
.INITVAL_36({2'b00, INIT[879*18 +: 18], 2'b00, INIT[878*18 +: 18], 2'b00, INIT[877*18 +: 18], 2'b00, INIT[876*18 +: 18], 
          2'b00, INIT[875*18 +: 18], 2'b00, INIT[874*18 +: 18], 2'b00, INIT[873*18 +: 18], 2'b00, INIT[872*18 +: 18], 
          2'b00, INIT[871*18 +: 18], 2'b00, INIT[870*18 +: 18], 2'b00, INIT[869*18 +: 18], 2'b00, INIT[868*18 +: 18], 
          2'b00, INIT[867*18 +: 18], 2'b00, INIT[866*18 +: 18], 2'b00, INIT[865*18 +: 18], 2'b00, INIT[864*18 +: 18]}),
.INITVAL_37({2'b00, INIT[895*18 +: 18], 2'b00, INIT[894*18 +: 18], 2'b00, INIT[893*18 +: 18], 2'b00, INIT[892*18 +: 18], 
          2'b00, INIT[891*18 +: 18], 2'b00, INIT[890*18 +: 18], 2'b00, INIT[889*18 +: 18], 2'b00, INIT[888*18 +: 18], 
          2'b00, INIT[887*18 +: 18], 2'b00, INIT[886*18 +: 18], 2'b00, INIT[885*18 +: 18], 2'b00, INIT[884*18 +: 18], 
          2'b00, INIT[883*18 +: 18], 2'b00, INIT[882*18 +: 18], 2'b00, INIT[881*18 +: 18], 2'b00, INIT[880*18 +: 18]}),
.INITVAL_38({2'b00, INIT[911*18 +: 18], 2'b00, INIT[910*18 +: 18], 2'b00, INIT[909*18 +: 18], 2'b00, INIT[908*18 +: 18], 
          2'b00, INIT[907*18 +: 18], 2'b00, INIT[906*18 +: 18], 2'b00, INIT[905*18 +: 18], 2'b00, INIT[904*18 +: 18], 
          2'b00, INIT[903*18 +: 18], 2'b00, INIT[902*18 +: 18], 2'b00, INIT[901*18 +: 18], 2'b00, INIT[900*18 +: 18], 
          2'b00, INIT[899*18 +: 18], 2'b00, INIT[898*18 +: 18], 2'b00, INIT[897*18 +: 18], 2'b00, INIT[896*18 +: 18]}),
.INITVAL_39({2'b00, INIT[927*18 +: 18], 2'b00, INIT[926*18 +: 18], 2'b00, INIT[925*18 +: 18], 2'b00, INIT[924*18 +: 18], 
          2'b00, INIT[923*18 +: 18], 2'b00, INIT[922*18 +: 18], 2'b00, INIT[921*18 +: 18], 2'b00, INIT[920*18 +: 18], 
          2'b00, INIT[919*18 +: 18], 2'b00, INIT[918*18 +: 18], 2'b00, INIT[917*18 +: 18], 2'b00, INIT[916*18 +: 18], 
          2'b00, INIT[915*18 +: 18], 2'b00, INIT[914*18 +: 18], 2'b00, INIT[913*18 +: 18], 2'b00, INIT[912*18 +: 18]}),
.INITVAL_3A({2'b00, INIT[943*18 +: 18], 2'b00, INIT[942*18 +: 18], 2'b00, INIT[941*18 +: 18], 2'b00, INIT[940*18 +: 18], 
          2'b00, INIT[939*18 +: 18], 2'b00, INIT[938*18 +: 18], 2'b00, INIT[937*18 +: 18], 2'b00, INIT[936*18 +: 18], 
          2'b00, INIT[935*18 +: 18], 2'b00, INIT[934*18 +: 18], 2'b00, INIT[933*18 +: 18], 2'b00, INIT[932*18 +: 18], 
          2'b00, INIT[931*18 +: 18], 2'b00, INIT[930*18 +: 18], 2'b00, INIT[929*18 +: 18], 2'b00, INIT[928*18 +: 18]}),
.INITVAL_3B({2'b00, INIT[959*18 +: 18], 2'b00, INIT[958*18 +: 18], 2'b00, INIT[957*18 +: 18], 2'b00, INIT[956*18 +: 18], 
          2'b00, INIT[955*18 +: 18], 2'b00, INIT[954*18 +: 18], 2'b00, INIT[953*18 +: 18], 2'b00, INIT[952*18 +: 18], 
          2'b00, INIT[951*18 +: 18], 2'b00, INIT[950*18 +: 18], 2'b00, INIT[949*18 +: 18], 2'b00, INIT[948*18 +: 18], 
          2'b00, INIT[947*18 +: 18], 2'b00, INIT[946*18 +: 18], 2'b00, INIT[945*18 +: 18], 2'b00, INIT[944*18 +: 18]}),
.INITVAL_3C({2'b00, INIT[975*18 +: 18], 2'b00, INIT[974*18 +: 18], 2'b00, INIT[973*18 +: 18], 2'b00, INIT[972*18 +: 18], 
          2'b00, INIT[971*18 +: 18], 2'b00, INIT[970*18 +: 18], 2'b00, INIT[969*18 +: 18], 2'b00, INIT[968*18 +: 18], 
          2'b00, INIT[967*18 +: 18], 2'b00, INIT[966*18 +: 18], 2'b00, INIT[965*18 +: 18], 2'b00, INIT[964*18 +: 18], 
          2'b00, INIT[963*18 +: 18], 2'b00, INIT[962*18 +: 18], 2'b00, INIT[961*18 +: 18], 2'b00, INIT[960*18 +: 18]}),
.INITVAL_3D({2'b00, INIT[991*18 +: 18], 2'b00, INIT[990*18 +: 18], 2'b00, INIT[989*18 +: 18], 2'b00, INIT[988*18 +: 18], 
          2'b00, INIT[987*18 +: 18], 2'b00, INIT[986*18 +: 18], 2'b00, INIT[985*18 +: 18], 2'b00, INIT[984*18 +: 18], 
          2'b00, INIT[983*18 +: 18], 2'b00, INIT[982*18 +: 18], 2'b00, INIT[981*18 +: 18], 2'b00, INIT[980*18 +: 18], 
          2'b00, INIT[979*18 +: 18], 2'b00, INIT[978*18 +: 18], 2'b00, INIT[977*18 +: 18], 2'b00, INIT[976*18 +: 18]}),
.INITVAL_3E({2'b00, INIT[1007*18 +: 18], 2'b00, INIT[1006*18 +: 18], 2'b00, INIT[1005*18 +: 18], 2'b00, INIT[1004*18 +: 18], 
          2'b00, INIT[1003*18 +: 18], 2'b00, INIT[1002*18 +: 18], 2'b00, INIT[1001*18 +: 18], 2'b00, INIT[1000*18 +: 18], 
          2'b00, INIT[999*18 +: 18], 2'b00, INIT[998*18 +: 18], 2'b00, INIT[997*18 +: 18], 2'b00, INIT[996*18 +: 18], 
          2'b00, INIT[995*18 +: 18], 2'b00, INIT[994*18 +: 18], 2'b00, INIT[993*18 +: 18], 2'b00, INIT[992*18 +: 18]}),
.INITVAL_3F({2'b00, INIT[1023*18 +: 18], 2'b00, INIT[1022*18 +: 18], 2'b00, INIT[1021*18 +: 18], 2'b00, INIT[1020*18 +: 18], 
          2'b00, INIT[1019*18 +: 18], 2'b00, INIT[1018*18 +: 18], 2'b00, INIT[1017*18 +: 18], 2'b00, INIT[1016*18 +: 18], 
          2'b00, INIT[1015*18 +: 18], 2'b00, INIT[1014*18 +: 18], 2'b00, INIT[1013*18 +: 18], 2'b00, INIT[1012*18 +: 18], 
          2'b00, INIT[1011*18 +: 18], 2'b00, INIT[1010*18 +: 18], 2'b00, INIT[1009*18 +: 18], 2'b00, INIT[1008*18 +: 18]}),
