    .ADA0(A1EN[0]), .ADA1(A1EN[1]), .ADA2(1'b0), .ADA3(1'b0), .ADA4(A1ADDR[0]), .ADA5(A1ADDR[1]), .ADA6(A1ADDR[2]), .ADA7(A1ADDR[3]), .ADA8(A1ADDR[4]), .ADA9(A1ADDR[5]), .ADA10(A1ADDR[6]), .ADA11(A1ADDR[7]), .ADA12(A1ADDR[8]), .ADA13(A1ADDR[9]),
    .ADB0(1'b0), .ADB1(1'b0), .ADB2(1'b0), .ADB3(1'b0), .ADB4(B1ADDR[0]), .ADB5(B1ADDR[1]), .ADB6(B1ADDR[2]), .ADB7(B1ADDR[3]), .ADB8(B1ADDR[4]), .ADB9(B1ADDR[5]), .ADB10(B1ADDR[6]), .ADB11(B1ADDR[7]), .ADB12(B1ADDR[8]), .ADB13(B1ADDR[9]),
    .DIA0(A1DATA[0]), .DIA1(A1DATA[1]), .DIA2(A1DATA[2]), .DIA3(A1DATA[3]), .DIA4(A1DATA[4]), .DIA5(A1DATA[5]), .DIA6(A1DATA[6]), .DIA7(A1DATA[7]), .DIA8(A1DATA[8]), .DIA9(A1DATA[9]), .DIA10(A1DATA[10]), .DIA11(A1DATA[11]), .DIA12(A1DATA[12]), .DIA13(A1DATA[13]), .DIA14(A1DATA[14]), .DIA15(A1DATA[15]), .DIA16(A1DATA[16]), .DIA17(A1DATA[17]),
    .DOB0(B1DATA[0]), .DOB1(B1DATA[1]), .DOB2(B1DATA[2]), .DOB3(B1DATA[3]), .DOB4(B1DATA[4]), .DOB5(B1DATA[5]), .DOB6(B1DATA[6]), .DOB7(B1DATA[7]), .DOB8(B1DATA[8]), .DOB9(B1DATA[9]), .DOB10(B1DATA[10]), .DOB11(B1DATA[11]), .DOB12(B1DATA[12]), .DOB13(B1DATA[13]), .DOB14(B1DATA[14]), .DOB15(B1DATA[15]), .DOB16(B1DATA[16]), .DOB17(B1DATA[17]),
